`define CYCLE_TIME 20

module PATTERN(
    // Output signals
    clk,
	rst_n,
	in_valid,
    in_xp_real, 
    in_xp_img,
    // Input signals
    out_valid, 
	out_yp_real,
    out_yp_img
);
// ========================================
// Input & Output
// ========================================
output reg clk, rst_n, in_valid;
output reg signed [15:0] in_xp_real, in_xp_img;

input out_valid;
input signed [15:0] out_yp_real, out_yp_img;

//================================================================
// clock
//================================================================
integer CYCLE;
initial begin 
    CYCLE = `CYCLE_TIME;
    clk = 0 ;
end
always #(`CYCLE_TIME/2.0) clk = ~clk;
//================================================================
// integer
//================================================================
integer pat_num, pat_tot;
integer latency;
integer total_latency = 0;
integer i, f_in, m;
integer a;

reg signed [15:0] STG_R [0:8][0:255];  // 9 個 stage (0~8)，每個 256 點
reg signed [15:0] STG_I [0:8][0:255];

reg[9:0] out_counter;
reg signed [15:0] xp_real_reg[0:255], xp_img_reg[0:255];
reg signed [15:0] golden_out_yp_img[0:255], golden_out_yp_real[0:255];

reg signed [15:0] in_real, in_img;

reg signed [15:0] w_real[0:255];
reg signed [15:0] w_img [0:255];

reg [8:0] idx[0:255];
/*
wire signed [31:0] xq_w_real0;
wire signed [31:0] xq_w_real1;
wire signed [31:0] xq_w_imag0;
wire signed [31:0] xq_w_imag1;
wire signed [31:0] xq_w_real ;
wire signed [31:0] xq_w_imag ;
wire signed [31:0] xp_real_scaled;
wire signed [31:0] xp_img_scaled;
wire signed [31:0] yp_real_scaled;
wire signed [31:0] yp_img_scaled ;
wire signed [31:0] yq_real_scaled;
wire signed [31:0] yq_img_scaled ;
*/
initial begin
    w_real[0] = 16'h7fff; // 1.0000
    w_img[0] = 16'h0000; // -0.0000
    w_real[1] = 16'h7ff6; // 0.9997
    w_img[1] = 16'hfcdc; // -0.0245
    w_real[2] = 16'h7fd9; // 0.9988
    w_img[2] = 16'hf9b8; // -0.0491
    w_real[3] = 16'h7fa7; // 0.9973
    w_img[3] = 16'hf695; // -0.0736
    w_real[4] = 16'h7f62; // 0.9952
    w_img[4] = 16'hf374; // -0.0980
    w_real[5] = 16'h7f0a; // 0.9925
    w_img[5] = 16'hf055; // -0.1224
    w_real[6] = 16'h7e9d; // 0.9892
    w_img[6] = 16'hed38; // -0.1467
    w_real[7] = 16'h7e1e; // 0.9853
    w_img[7] = 16'hea1e; // -0.1710
    w_real[8] = 16'h7d8a; // 0.9808
    w_img[8] = 16'he707; // -0.1951
    w_real[9] = 16'h7ce4; // 0.9757
    w_img[9] = 16'he3f4; // -0.2191
    w_real[10] = 16'h7c2a; // 0.9700
    w_img[10] = 16'he0e6; // -0.2430
    w_real[11] = 16'h7b5d; // 0.9638
    w_img[11] = 16'hdddc; // -0.2667
    w_real[12] = 16'h7a7d; // 0.9569
    w_img[12] = 16'hdad8; // -0.2903
    w_real[13] = 16'h798a; // 0.9495
    w_img[13] = 16'hd7d9; // -0.3137
    w_real[14] = 16'h7885; // 0.9415
    w_img[14] = 16'hd4e1; // -0.3369
    w_real[15] = 16'h776c; // 0.9330
    w_img[15] = 16'hd1ef; // -0.3599
    w_real[16] = 16'h7642; // 0.9239
    w_img[16] = 16'hcf04; // -0.3827
    w_real[17] = 16'h7505; // 0.9142
    w_img[17] = 16'hcc21; // -0.4052
    w_real[18] = 16'h73b6; // 0.9040
    w_img[18] = 16'hc946; // -0.4276
    w_real[19] = 16'h7255; // 0.8932
    w_img[19] = 16'hc673; // -0.4496
    w_real[20] = 16'h70e3; // 0.8819
    w_img[20] = 16'hc3a9; // -0.4714
    w_real[21] = 16'h6f5f; // 0.8701
    w_img[21] = 16'hc0e9; // -0.4929
    w_real[22] = 16'h6dca; // 0.8577
    w_img[22] = 16'hbe32; // -0.5141
    w_real[23] = 16'h6c24; // 0.8449
    w_img[23] = 16'hbb85; // -0.5350
    w_real[24] = 16'h6a6e; // 0.8315
    w_img[24] = 16'hb8e3; // -0.5556
    w_real[25] = 16'h68a7; // 0.8176
    w_img[25] = 16'hb64c; // -0.5758
    w_real[26] = 16'h66d0; // 0.8032
    w_img[26] = 16'hb3c0; // -0.5957
    w_real[27] = 16'h64e9; // 0.7883
    w_img[27] = 16'hb140; // -0.6152
    w_real[28] = 16'h62f2; // 0.7730
    w_img[28] = 16'haecc; // -0.6344
    w_real[29] = 16'h60ec; // 0.7572
    w_img[29] = 16'hac65; // -0.6532
    w_real[30] = 16'h5ed7; // 0.7410
    w_img[30] = 16'haa0a; // -0.6716
    w_real[31] = 16'h5cb4; // 0.7242
    w_img[31] = 16'ha7bd; // -0.6895
    w_real[32] = 16'h5a82; // 0.7071
    w_img[32] = 16'ha57e; // -0.7071
    w_real[33] = 16'h5843; // 0.6895
    w_img[33] = 16'ha34c; // -0.7242
    w_real[34] = 16'h55f6; // 0.6716
    w_img[34] = 16'ha129; // -0.7410
    w_real[35] = 16'h539b; // 0.6532
    w_img[35] = 16'h9f14; // -0.7572
    w_real[36] = 16'h5134; // 0.6344
    w_img[36] = 16'h9d0e; // -0.7730
    w_real[37] = 16'h4ec0; // 0.6152
    w_img[37] = 16'h9b17; // -0.7883
    w_real[38] = 16'h4c40; // 0.5957
    w_img[38] = 16'h9930; // -0.8032
    w_real[39] = 16'h49b4; // 0.5758
    w_img[39] = 16'h9759; // -0.8176
    w_real[40] = 16'h471d; // 0.5556
    w_img[40] = 16'h9592; // -0.8315
    w_real[41] = 16'h447b; // 0.5350
    w_img[41] = 16'h93dc; // -0.8449
    w_real[42] = 16'h41ce; // 0.5141
    w_img[42] = 16'h9236; // -0.8577
    w_real[43] = 16'h3f17; // 0.4929
    w_img[43] = 16'h90a1; // -0.8701
    w_real[44] = 16'h3c57; // 0.4714
    w_img[44] = 16'h8f1d; // -0.8819
    w_real[45] = 16'h398d; // 0.4496
    w_img[45] = 16'h8dab; // -0.8932
    w_real[46] = 16'h36ba; // 0.4276
    w_img[46] = 16'h8c4a; // -0.9040
    w_real[47] = 16'h33df; // 0.4052
    w_img[47] = 16'h8afb; // -0.9142
    w_real[48] = 16'h30fc; // 0.3827
    w_img[48] = 16'h89be; // -0.9239
    w_real[49] = 16'h2e11; // 0.3599
    w_img[49] = 16'h8894; // -0.9330
    w_real[50] = 16'h2b1f; // 0.3369
    w_img[50] = 16'h877b; // -0.9415
    w_real[51] = 16'h2827; // 0.3137
    w_img[51] = 16'h8676; // -0.9495
    w_real[52] = 16'h2528; // 0.2903
    w_img[52] = 16'h8583; // -0.9569
    w_real[53] = 16'h2224; // 0.2667
    w_img[53] = 16'h84a3; // -0.9638
    w_real[54] = 16'h1f1a; // 0.2430
    w_img[54] = 16'h83d6; // -0.9700
    w_real[55] = 16'h1c0c; // 0.2191
    w_img[55] = 16'h831c; // -0.9757
    w_real[56] = 16'h18f9; // 0.1951
    w_img[56] = 16'h8276; // -0.9808
    w_real[57] = 16'h15e2; // 0.1710
    w_img[57] = 16'h81e2; // -0.9853
    w_real[58] = 16'h12c8; // 0.1467
    w_img[58] = 16'h8163; // -0.9892
    w_real[59] = 16'h0fab; // 0.1224
    w_img[59] = 16'h80f6; // -0.9925
    w_real[60] = 16'h0c8c; // 0.0980
    w_img[60] = 16'h809e; // -0.9952
    w_real[61] = 16'h096b; // 0.0736
    w_img[61] = 16'h8059; // -0.9973
    w_real[62] = 16'h0648; // 0.0491
    w_img[62] = 16'h8027; // -0.9988
    w_real[63] = 16'h0324; // 0.0245
    w_img[63] = 16'h800a; // -0.9997
    w_real[64] = 16'h0000; // 0.0000
    w_img[64] = 16'h8000; // -1.0000
    w_real[65] = 16'hfcdc; // -0.0245
    w_img[65] = 16'h800a; // -0.9997
    w_real[66] = 16'hf9b8; // -0.0491
    w_img[66] = 16'h8027; // -0.9988
    w_real[67] = 16'hf695; // -0.0736
    w_img[67] = 16'h8059; // -0.9973
    w_real[68] = 16'hf374; // -0.0980
    w_img[68] = 16'h809e; // -0.9952
    w_real[69] = 16'hf055; // -0.1224
    w_img[69] = 16'h80f6; // -0.9925
    w_real[70] = 16'hed38; // -0.1467
    w_img[70] = 16'h8163; // -0.9892
    w_real[71] = 16'hea1e; // -0.1710
    w_img[71] = 16'h81e2; // -0.9853
    w_real[72] = 16'he707; // -0.1951
    w_img[72] = 16'h8276; // -0.9808
    w_real[73] = 16'he3f4; // -0.2191
    w_img[73] = 16'h831c; // -0.9757
    w_real[74] = 16'he0e6; // -0.2430
    w_img[74] = 16'h83d6; // -0.9700
    w_real[75] = 16'hdddc; // -0.2667
    w_img[75] = 16'h84a3; // -0.9638
    w_real[76] = 16'hdad8; // -0.2903
    w_img[76] = 16'h8583; // -0.9569
    w_real[77] = 16'hd7d9; // -0.3137
    w_img[77] = 16'h8676; // -0.9495
    w_real[78] = 16'hd4e1; // -0.3369
    w_img[78] = 16'h877b; // -0.9415
    w_real[79] = 16'hd1ef; // -0.3599
    w_img[79] = 16'h8894; // -0.9330
    w_real[80] = 16'hcf04; // -0.3827
    w_img[80] = 16'h89be; // -0.9239
    w_real[81] = 16'hcc21; // -0.4052
    w_img[81] = 16'h8afb; // -0.9142
    w_real[82] = 16'hc946; // -0.4276
    w_img[82] = 16'h8c4a; // -0.9040
    w_real[83] = 16'hc673; // -0.4496
    w_img[83] = 16'h8dab; // -0.8932
    w_real[84] = 16'hc3a9; // -0.4714
    w_img[84] = 16'h8f1d; // -0.8819
    w_real[85] = 16'hc0e9; // -0.4929
    w_img[85] = 16'h90a1; // -0.8701
    w_real[86] = 16'hbe32; // -0.5141
    w_img[86] = 16'h9236; // -0.8577
    w_real[87] = 16'hbb85; // -0.5350
    w_img[87] = 16'h93dc; // -0.8449
    w_real[88] = 16'hb8e3; // -0.5556
    w_img[88] = 16'h9592; // -0.8315
    w_real[89] = 16'hb64c; // -0.5758
    w_img[89] = 16'h9759; // -0.8176
    w_real[90] = 16'hb3c0; // -0.5957
    w_img[90] = 16'h9930; // -0.8032
    w_real[91] = 16'hb140; // -0.6152
    w_img[91] = 16'h9b17; // -0.7883
    w_real[92] = 16'haecc; // -0.6344
    w_img[92] = 16'h9d0e; // -0.7730
    w_real[93] = 16'hac65; // -0.6532
    w_img[93] = 16'h9f14; // -0.7572
    w_real[94] = 16'haa0a; // -0.6716
    w_img[94] = 16'ha129; // -0.7410
    w_real[95] = 16'ha7bd; // -0.6895
    w_img[95] = 16'ha34c; // -0.7242
    w_real[96] = 16'ha57e; // -0.7071
    w_img[96] = 16'ha57e; // -0.7071
    w_real[97] = 16'ha34c; // -0.7242
    w_img[97] = 16'ha7bd; // -0.6895
    w_real[98] = 16'ha129; // -0.7410
    w_img[98] = 16'haa0a; // -0.6716
    w_real[99] = 16'h9f14; // -0.7572
    w_img[99] = 16'hac65; // -0.6532
    w_real[100] = 16'h9d0e; // -0.7730
    w_img[100] = 16'haecc; // -0.6344
    w_real[101] = 16'h9b17; // -0.7883
    w_img[101] = 16'hb140; // -0.6152
    w_real[102] = 16'h9930; // -0.8032
    w_img[102] = 16'hb3c0; // -0.5957
    w_real[103] = 16'h9759; // -0.8176
    w_img[103] = 16'hb64c; // -0.5758
    w_real[104] = 16'h9592; // -0.8315
    w_img[104] = 16'hb8e3; // -0.5556
    w_real[105] = 16'h93dc; // -0.8449
    w_img[105] = 16'hbb85; // -0.5350
    w_real[106] = 16'h9236; // -0.8577
    w_img[106] = 16'hbe32; // -0.5141
    w_real[107] = 16'h90a1; // -0.8701
    w_img[107] = 16'hc0e9; // -0.4929
    w_real[108] = 16'h8f1d; // -0.8819
    w_img[108] = 16'hc3a9; // -0.4714
    w_real[109] = 16'h8dab; // -0.8932
    w_img[109] = 16'hc673; // -0.4496
    w_real[110] = 16'h8c4a; // -0.9040
    w_img[110] = 16'hc946; // -0.4276
    w_real[111] = 16'h8afb; // -0.9142
    w_img[111] = 16'hcc21; // -0.4052
    w_real[112] = 16'h89be; // -0.9239
    w_img[112] = 16'hcf04; // -0.3827
    w_real[113] = 16'h8894; // -0.9330
    w_img[113] = 16'hd1ef; // -0.3599
    w_real[114] = 16'h877b; // -0.9415
    w_img[114] = 16'hd4e1; // -0.3369
    w_real[115] = 16'h8676; // -0.9495
    w_img[115] = 16'hd7d9; // -0.3137
    w_real[116] = 16'h8583; // -0.9569
    w_img[116] = 16'hdad8; // -0.2903
    w_real[117] = 16'h84a3; // -0.9638
    w_img[117] = 16'hdddc; // -0.2667
    w_real[118] = 16'h83d6; // -0.9700
    w_img[118] = 16'he0e6; // -0.2430
    w_real[119] = 16'h831c; // -0.9757
    w_img[119] = 16'he3f4; // -0.2191
    w_real[120] = 16'h8276; // -0.9808
    w_img[120] = 16'he707; // -0.1951
    w_real[121] = 16'h81e2; // -0.9853
    w_img[121] = 16'hea1e; // -0.1710
    w_real[122] = 16'h8163; // -0.9892
    w_img[122] = 16'hed38; // -0.1467
    w_real[123] = 16'h80f6; // -0.9925
    w_img[123] = 16'hf055; // -0.1224
    w_real[124] = 16'h809e; // -0.9952
    w_img[124] = 16'hf374; // -0.0980
    w_real[125] = 16'h8059; // -0.9973
    w_img[125] = 16'hf695; // -0.0736
    w_real[126] = 16'h8027; // -0.9988
    w_img[126] = 16'hf9b8; // -0.0491
    w_real[127] = 16'h800a; // -0.9997
    w_img[127] = 16'hfcdc; // -0.0245    
    for (m = 0; m < 128; m = m + 1) begin
        w_real[m+128] = -w_real[m];
        w_img[m+128]  = -w_img[m];
    end    
end
initial begin
    // Initialize signals
    reset_task;
    pat_tot = 10000;
    for (i = 0 ; i < 256; i = i+1) begin
        xp_real_reg[i] = 0;
        xp_img_reg[i] = 0;
    end
    
    for(pat_num = 0; pat_num < pat_tot; pat_num = pat_num + 1) begin
        input_task;
        @(negedge clk);
        in_valid = 1;
        for (i = 0 ; i < 256 ; i = i + 1 ) begin
            in_xp_real = xp_real_reg[i];
            in_xp_img = xp_img_reg[i];
            @(negedge clk);
        end
        @(negedge clk);
        in_valid = 0;
        in_xp_real = 'bx;
        in_xp_img = 'bx;
        latency = 0;

        conjugate_task;
        cal_gold_task;
        wait_out_valid_task;
        check_ans_task;
        $display("\033[0;34mPASS SET NO.%4d,\033[m \033[0;32m     Execution Cycle: %3d\033[m", pat_num, latency);
    end
	display_pass;
	$finish;
end
localparam integer SHIFT = 15;  // 要跟 RTL module 的 parameter 一致

task automatic butterfly(
    input  signed [15:0] xp_real,
    input  signed [15:0] xp_img,
    input  signed [15:0] xq_real,
    input  signed [15:0] xq_img,
    input  signed [15:0] w_real,
    input  signed [15:0] w_img,
    output signed [15:0] yp_real,
    output signed [15:0] yp_img,
    output signed [15:0] yq_real,
    output signed [15:0] yq_img
);
    integer xq_w_r0, xq_w_r1, xq_w_i0, xq_w_i1;
    integer xq_w_r,  xq_w_i;
    integer xp_r_scaled, xp_i_scaled;
    integer yp_r_scaled, yp_i_scaled;
    integer yq_r_scaled, yq_i_scaled;
    integer tmp;
begin
    // 1) xq * W  (跟 RTL 一樣)
    xq_w_r0 = xq_real * w_real;
    xq_w_r1 = xq_img  * w_img;
    xq_w_i0 = xq_real * w_img;
    xq_w_i1 = xq_img  * w_real;

    xq_w_r  = xq_w_r0 - xq_w_r1;
    xq_w_i  = xq_w_i0 + xq_w_i1;

    // 2) xp 先 sign-extend 再 shift，模仿 RTL
    xp_r_scaled = $signed({{16{xp_real[15]}}, xp_real}) <<< SHIFT;
    xp_i_scaled = $signed({{16{xp_img[15]}},  xp_img }) <<< SHIFT;

    // 3) butterfly
    yp_r_scaled = xp_r_scaled + xq_w_r;
    yp_i_scaled = xp_i_scaled + xq_w_i;
    yq_r_scaled = xp_r_scaled - xq_w_r;
    yq_i_scaled = xp_i_scaled - xq_w_i;

    // 4) >> SHIFT 再取 16-bit（跟 RTL 的 [SHIFT+15:SHIFT] 等價）
    tmp     = yp_r_scaled >>> SHIFT;
    yp_real = tmp[15:0];

    tmp     = yp_i_scaled >>> SHIFT;
    yp_img  = tmp[15:0];

    tmp     = yq_r_scaled >>> SHIFT;
    yq_real = tmp[15:0];

    tmp     = yq_i_scaled >>> SHIFT;
    yq_img  = tmp[15:0];
end
endtask

function integer bitrev8(input integer x);
    integer i;
    integer r;
begin
    r = 0;
    for (i = 0; i < 8; i = i + 1) begin
        r = r | (((x >> i) & 1) << (7 - i));
    end
    bitrev8 = r;
end
endfunction

task cal_gold_task; begin
    fft_task;
    for (i = 0 ; i < 256; i = i + 1) begin
            golden_out_yp_real[n] = (temp_golden_out_yp_real[n])/256;
            golden_out_yp_img[n]  = (-temp_golden_out_yp_img[n])/256; 
    end
end
endtask

task fft_task;
    integer N;
    integer STAGES;
    integer s, n, g, j;
    integer dista, group_size, num_groups;
    integer p, q, tw_idx;
    reg signed [15:0] xp_r, xp_i, xq_r, xq_i;
    reg signed [15:0] w_r, w_i;
    integer bits, b, g_br;
begin
    N       = 256;
    STAGES  = 8;

    // 0) stage0 接 DUT 的 input
    for (n = 0; n < N; n = n + 1) begin
        STG_R[0][n] = xp_real_reg[n];  // Q1.15
        STG_I[0][n] = -xp_img_reg[n];
    end

    // 1) 8 個 stage，DIF + 你的 wiring + twiddle 排法
    for (s = 0; s < STAGES; s = s + 1) begin
        // 每層距離: 第一層 128, 第二層 64, ..., 第八層 1
        dista = N >> (s + 1);       // 128,64,32,16,8,4,2,1
        group_size  = dista << 1;          // 256,128,64,32,16,8,4,2
        num_groups  = N / group_size;     // 1,2,4,8,16,32,64,128

        bits = s; // 用 s 個 bits 來做 group index 的 bit-reverse

        for (g = 0; g < num_groups; g = g + 1) begin
            // ---- group twiddle index ----
            g_br = 0;
            for (b = 0; b < bits; b = b + 1) begin
                g_br = g_br | (((g >> b) & 1) << (bits - 1 - b));
            end
            // stage0 (s=0) 時 bits=0 → g_br=0 → tw_idx=0 → 全部 w[0]
            tw_idx = g_br * dista;  // stage1: dist=64, g=0,1 → 0,64
            w_r    = w_real[tw_idx];
            w_i    = w_img [tw_idx];

            // ---- 這個 group 裡的 dist 個 butterfly ----
            for (j = 0; j < dista; j = j + 1) begin
                p = g * group_size + j;
                q = p + dista;

                xp_r = STG_R[s][p];
                xp_i = STG_I[s][p];
                xq_r = STG_R[s][q];
                xq_i = STG_I[s][q];
                /*
                if (s==0 && g==0 && j==0) begin
                    $display("GOLDEN stage0 first butterfly:");
                    $display("xp_r=%h xp_i=%h", xp_r, xp_i);
                    $display("xq_r=%h xq_i=%h", xq_r, xq_i);
                    $display("dist=%0d tw_idx=%0d w_r=%h w_i=%h", dista, tw_idx, w_r, w_i);
                end
                */
                butterfly(
                    xp_r, xp_i,
                    xq_r, xq_i,
                    w_r,  w_i,
                    STG_R[s+1][p], STG_I[s+1][p],
                    STG_R[s+1][q], STG_I[s+1][q]
                );
                /*
                if (s==0 && g==0 && j==0) begin
                    $display("golden yp_r=%h yp_i=%h", STG_R[1][0], STG_I[1][0]);
                end
                */
            end
        end
    end

    // 2) 輸出 stage 8 的結果（假設 DUT 也是 bit-reversed order）
    for (n = 0; n < N; n = n + 1) begin
        temp_golden_out_yp_real[n] = STG_R[STAGES][bitrev8(n)][15:0];
        temp_golden_out_yp_img[n]  = STG_I[STAGES][bitrev8(n)][15:0];
    end
end
endtask


task check_ans_task; begin
    
    out_counter = 0;
    while(out_valid !== 1'b0) begin
        if(out_yp_real !== golden_out_yp_real[out_counter]) begin
            $display("***************************************************************************");
            $display("                         Your answer is incorrect! (real)                        ");
            $display("                         failed at cycle = %4d                         ", out_counter);
            $display("     Your answer = %4h", out_yp_real, "     Golden answer = %4h", golden_out_yp_real[out_counter]);
            $display("***************************************************************************");
            $finish;
        end
        else if(out_yp_img !== golden_out_yp_img[out_counter]) begin
            $display("***************************************************************************");
            $display("                         Your answer is incorrect! (img)                         ");
            $display("                         failed at cycle = %4d                         ", out_counter);
            $display("     Your answer = %4h", out_yp_img, "     Golden answer = %4h", golden_out_yp_img[out_counter]);
            $display("***************************************************************************");
            $finish;
        end

        @(negedge clk);
        out_counter = out_counter + 1;
    end
    if (out_counter != 256) begin
        $display("***************************************************************************");
        $display("            Your out_valid should be pulled up for 256 cycles!             ");
        $display("     Your answer = %4d", out_counter, "     Golden answer = 256");
        $display("***************************************************************************");
        $finish;
    end
end
endtask



task wait_out_valid_task; begin
    latency =0;
    while (out_valid === 0) begin
        latency = latency + 1;
        if (latency == (1000*CYCLE)) begin // max latency = 1000
            $display("                    OVER 1000 LATENCY                   ");
            repeat (2) @(negedge clk);
            $finish;
        end
        @(negedge clk);
    end
    total_latency = total_latency + latency;
end 
endtask

task input_task; begin
    
    for (i = 0 ; i < 256 ; i = i + 1) begin
        xp_real_reg[i] = $urandom_range(-32768, 32767);
        xp_img_reg[i] = $urandom_range(-32768, 32767);
    end
    
    /*
    f_in  = $fopen("fft_input_q15_hex.txt", "r");
    if (f_in == 0) begin
        $display("Failed to open input.txt");
        $finish;
    end
    // Initialize signals

    for(i = 0 ; i < 256 ; i = i + 1)begin
        a = $fscanf(f_in, "%h %h", in_real, in_img);
		xp_real_reg[i] = in_real;
		xp_img_reg[i] = in_img;
    end
    */
end
endtask

task reset_task;begin
    rst_n = 1'b1;
    in_valid = 1'b0;
	in_xp_real = 16'bx;
    in_xp_img = 16'bx;
    total_latency = 0;

    // Apply reset
    #CYCLE; rst_n = 1'b0; 
    #CYCLE; rst_n = 1'b1;
	#(100-CYCLE); 

	//@(negedge clk);   
    // Check initial conditions
    if (out_valid !== 1'b0 || out_yp_img !== 16'b00000000 || out_yp_real !== 16'b0000) begin
        $display("                    RESET TASK FAIL                   ");
        repeat (2) #CYCLE;
        $finish;
    end
    #CYCLE; 

	
end
endtask

task display_pass; begin
	$display("[38;2;178;138;79m&[0m[38;2;179;139;79m&[0m[38;2;179;139;80m&[0m[38;2;180;140;80m&[0m[38;2;180;140;80m&[0m[38;2;180;140;81m&[0m[38;2;180;140;81m&[0m[38;2;181;141;82m&[0m[38;2;181;141;82m&[0m[38;2;181;141;81m&[0m[38;2;183;143;82m&[0m[38;2;183;143;83m&[0m[38;2;182;142;82m&[0m[38;2;182;142;82m&[0m[38;2;183;143;83m&[0m[38;2;184;144;84m&[0m[38;2;184;144;82m&[0m[38;2;183;143;81m&[0m[38;2;183;143;83m&[0m[38;2;183;143;84m&[0m[38;2;183;143;84m&[0m[38;2;183;143;84m&[0m[38;2;184;144;85m&[0m[38;2;183;143;84m&[0m[38;2;183;143;84m&[0m[38;2;183;143;84m&[0m[38;2;184;144;85m&[0m[38;2;184;144;85m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;183;143;82m&[0m[38;2;183;143;82m&[0m[38;2;184;144;83m&[0m[38;2;183;143;82m&[0m[38;2;183;143;83m&[0m[38;2;181;142;79m&[0m[38;2;181;137;78m&[0m[38;2;116;60;35mH[0m[38;2;75;7;6mX[0m[38;2;77;7;9mX[0m[38;2;70;9;7mX[0m[38;2;67;22;11mA[0m[38;2;89;60;41mM[0m[38;2;124;104;78m9[0m[38;2;169;150;116m@[0m[38;2;190;172;134m@[0m[38;2;192;174;136m@[0m[38;2;192;176;138m@[0m[38;2;192;177;136m@[0m[38;2;194;179;136m@[0m[38;2;201;186;146m@[0m[38;2;180;164;127m@[0m[38;2;186;170;134m@[0m[38;2;192;177;139m@[0m[38;2;196;181;142m@[0m[38;2;195;180;140m@[0m[38;2;196;181;141m@[0m[38;2;195;180;141m@[0m[38;2;195;180;141m@[0m[38;2;196;181;142m@[0m[38;2;194;179;140m@[0m[38;2;196;179;139m@[0m[38;2;196;178;138m@[0m[38;2;188;170;132m@[0m[38;2;164;145;112m&[0m[38;2;135;115;87mB[0m[38;2;94;74;52mH[0m[38;2;57;39;23m2[0m[38;2;47;22;13ms[0m[38;2;58;19;13mX[0m[38;2;74;17;13mA[0m[38;2;83;13;10mA[0m[38;2;91;12;11mA[0m[38;2;95;13;10m2[0m[38;2;92;14;9m2[0m[38;2;91;14;10m2[0m[38;2;89;10;12mA[0m[38;2;89;10;12mA[0m[38;2;85;14;6mA[0m[38;2;101;38;19m3[0m[38;2;148;93;61m9[0m[38;2;165;117;70mB[0m[38;2;159;117;63mB[0m[38;2;159;117;66mB[0m[38;2;159;118;66mB[0m[38;2;157;116;63mB[0m[38;2;156;115;64mB[0m[38;2;156;114;63mB[0m[38;2;157;115;65mB[0m[38;2;170;128;80m&[0m[38;2;171;129;81m&[0m[38;2;171;129;81m&[0m[38;2;172;130;82m&[0m[38;2;173;130;82m&[0m[38;2;148;111;66m9[0m[38;2;115;83;44mG[0m[38;2;135;94;56m#[0m[38;2;161;116;71mB[0m[38;2;177;137;87m&[0m[38;2;185;148;95m@[0m[38;2;187;152;95m@[0m[38;2;187;152;96m@[0m[38;2;188;151;96m@[0m[38;2;188;151;96m@[0m[38;2;188;151;96m@[0m[38;2;189;152;96m@[0m[38;2;187;150;95m@[0m[38;2;187;151;94m@[0m[38;2;187;151;92m@[0m[38;2;187;151;92m@[0m[38;2;188;151;96m@[0m[38;2;162;125;73mB[0m[38;2;143;104;57m9[0m[38;2;145;103;58m9[0m[38;2;146;103;59m9[0m[38;2;145;103;60m9[0m[38;2;143;100;58m9[0m[38;2;160;117;69mB[0m[38;2;177;138;79m&[0m[38;2;193;156;94m@[0m[38;2;194;157;99m@[0m[38;2;177;136;80m&[0m[38;2;183;141;87m&[0m[38;2;188;150;91m@[0m[38;2;186;152;87m&[0m[38;2;186;152;90m@[0m[38;2;185;149;87m&[0m");
	$display("[38;2;175;135;79m&[0m[38;2;176;136;80m&[0m[38;2;176;136;80m&[0m[38;2;177;137;81m&[0m[38;2;177;137;81m&[0m[38;2;177;138;80m&[0m[38;2;177;138;80m&[0m[38;2;178;138;81m&[0m[38;2;179;139;81m&[0m[38;2;178;139;80m&[0m[38;2;179;140;81m&[0m[38;2;180;140;82m&[0m[38;2;179;140;81m&[0m[38;2;179;140;81m&[0m[38;2;180;140;81m&[0m[38;2;181;141;81m&[0m[38;2;181;141;81m&[0m[38;2;181;141;80m&[0m[38;2;181;141;81m&[0m[38;2;181;141;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;82m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;181;141;80m&[0m[38;2;180;140;79m&[0m[38;2;181;141;80m&[0m[38;2;182;142;81m&[0m[38;2;181;140;79m&[0m[38;2;180;139;76m&[0m[38;2;181;140;77m&[0m[38;2;155;105;63m9[0m[38;2;81;17;8mA[0m[38;2;79;5;9mX[0m[38;2;71;4;4ms[0m[38;2;74;26;15m2[0m[38;2;125;97;72m#[0m[38;2;168;150;116m@[0m[38;2;182;164;127m@[0m[38;2;195;177;139m@[0m[38;2;186;168;130m@[0m[38;2;194;176;138m@[0m[38;2;192;175;139m@[0m[38;2;190;175;136m@[0m[38;2;208;193;154m@[0m[38;2;176;161;124m@[0m[38;2;181;165;131m@[0m[38;2;177;161;128m@[0m[38;2;190;175;138m@[0m[38;2;211;196;156m@[0m[38;2;195;180;142m@[0m[38;2;175;159;123m@[0m[38;2;189;174;136m@[0m[38;2;195;180;138m@[0m[38;2;201;186;146m@[0m[38;2;202;186;149m@[0m[38;2;193;177;138m@[0m[38;2;195;179;140m@[0m[38;2;204;188;150m@[0m[38;2;205;188;150m@[0m[38;2;189;173;134m@[0m[38;2;185;168;131m@[0m[38;2;167;151;116m@[0m[38;2;122;106;78m9[0m[38;2;77;57;38mh[0m[38;2;50;29;13mX[0m[38;2;50;20;9ms[0m[38;2;65;16;12mX[0m[38;2;78;12;10mA[0m[38;2;85;12;7mA[0m[38;2;84;11;5mA[0m[38;2;83;8;6mX[0m[38;2;83;8;9mA[0m[38;2;83;7;6mX[0m[38;2;82;8;5mX[0m[38;2;88;21;12m2[0m[38;2;132;76;48mS[0m[38;2;157;112;67mB[0m[38;2;155;115;64mB[0m[38;2;155;114;64mB[0m[38;2;155;113;64mB[0m[38;2;154;112;63m9[0m[38;2;153;111;63m9[0m[38;2;155;112;65mB[0m[38;2;170;128;80m&[0m[38;2;172;130;82m&[0m[38;2;173;131;83m&[0m[38;2;173;131;83m&[0m[38;2;174;131;84m&[0m[38;2;147;109;65m9[0m[38;2;113;80;42mG[0m[38;2;134;92;56m#[0m[38;2;160;115;71mB[0m[38;2;175;135;86m&[0m[38;2;186;149;96m@[0m[38;2;187;152;95m@[0m[38;2;186;151;94m@[0m[38;2;187;150;95m@[0m[38;2;186;151;96m@[0m[38;2;186;151;96m@[0m[38;2;186;151;96m@[0m[38;2;185;150;95m@[0m[38;2;186;149;94m@[0m[38;2;186;149;93m@[0m[38;2;186;149;93m@[0m[38;2;187;150;97m@[0m[38;2;162;125;74mB[0m[38;2;143;104;58m9[0m[38;2;145;103;58m9[0m[38;2;146;103;59m9[0m[38;2;145;103;60m9[0m[38;2;143;101;58m9[0m[38;2;155;113;66mB[0m[38;2;171;131;77m&[0m[38;2;186;149;91m&[0m[38;2;187;151;94m@[0m[38;2;167;128;74mB[0m[38;2;172;132;82m&[0m[38;2;183;144;92m&[0m[38;2;178;141;89m&[0m[38;2;150;113;72mB[0m[38;2;109;78;48mG[0m");
	$display("[38;2;173;134;80m&[0m[38;2;173;134;80m&[0m[38;2;173;134;80m&[0m[38;2;174;135;81m&[0m[38;2;174;135;80m&[0m[38;2;175;136;80m&[0m[38;2;176;137;81m&[0m[38;2;176;137;80m&[0m[38;2;176;138;80m&[0m[38;2;177;138;80m&[0m[38;2;177;138;81m&[0m[38;2;177;138;81m&[0m[38;2;177;138;81m&[0m[38;2;177;138;81m&[0m[38;2;178;137;81m&[0m[38;2;178;138;81m&[0m[38;2;178;138;81m&[0m[38;2;179;138;81m&[0m[38;2;179;139;81m&[0m[38;2;179;139;80m&[0m[38;2;179;139;80m&[0m[38;2;179;139;80m&[0m[38;2;179;139;80m&[0m[38;2;179;139;80m&[0m[38;2;180;140;80m&[0m[38;2;180;140;80m&[0m[38;2;180;140;80m&[0m[38;2;180;140;79m&[0m[38;2;180;140;79m&[0m[38;2;181;141;79m&[0m[38;2;180;140;79m&[0m[38;2;180;140;79m&[0m[38;2;180;140;79m&[0m[38;2;179;139;78m&[0m[38;2;179;139;78m&[0m[38;2;179;139;78m&[0m[38;2;180;140;79m&[0m[38;2;179;139;78m&[0m[38;2;179;139;78m&[0m[38;2;179;139;78m&[0m[38;2;178;138;77m&[0m[38;2;179;137;79m&[0m[38;2;178;137;77m&[0m[38;2;176;135;79m&[0m[38;2;122;66;41mG[0m[38;2;75;7;7mX[0m[38;2;70;2;3ms[0m[38;2;76;24;14mA[0m[38;2;162;130;105m&[0m[38;2;188;169;133m@[0m[38;2;168;152;112m@[0m[38;2;193;176;140m@[0m[38;2;183;167;130m@[0m[38;2;190;174;136m@[0m[38;2;192;176;137m@[0m[38;2;188;172;134m@[0m[38;2;208;192;157m@[0m[38;2;177;161;127m@[0m[38;2;145;129;94mB[0m[38;2;176;160;127m@[0m[38;2;178;163;129m@[0m[38;2;203;188;150m@[0m[38;2;216;199;160m@[0m[38;2;186;168;134m@[0m[38;2;123;105;74m9[0m[38;2;105;89;58mS[0m[38;2;183;168;132m@[0m[38;2;194;179;138m@[0m[38;2;211;195;160m@[0m[38;2;201;185;150m@[0m[38;2;171;155;120m@[0m[38;2;190;174;141m@[0m[38;2;205;189;153m@[0m[38;2;211;196;157m@[0m[38;2;192;176;135m@[0m[38;2;190;174;132m@[0m[38;2;196;180;139m@[0m[38;2;187;171;134m@[0m[38;2;154;139;107m&[0m[38;2;91;78;52mH[0m[38;2;47;31;15mX[0m[38;2;48;19;13ms[0m[38;2;59;14;13mX[0m[38;2;70;10;6mX[0m[38;2;76;7;5mX[0m[38;2;80;6;5mX[0m[38;2;81;8;6mX[0m[38;2;83;9;7mX[0m[38;2;81;7;4mX[0m[38;2;76;13;3mX[0m[38;2;120;70;46mG[0m[38;2;152;111;64m9[0m[38;2;153;112;61m9[0m[38;2;152;110;62m9[0m[38;2;152;110;62m9[0m[38;2;151;109;62m9[0m[38;2;153;110;64m9[0m[38;2;170;128;80m&[0m[38;2;173;131;83m&[0m[38;2;173;132;84m&[0m[38;2;173;132;84m&[0m[38;2;174;133;85m&[0m[38;2;146;109;66m9[0m[38;2;113;78;41mG[0m[38;2;131;92;55m#[0m[38;2;157;114;71mB[0m[38;2;174;133;84m&[0m[38;2;184;147;95m&[0m[38;2;185;151;95m@[0m[38;2;183;150;94m&[0m[38;2;185;149;96m@[0m[38;2;184;150;96m@[0m[38;2;184;150;96m@[0m[38;2;184;150;96m@[0m[38;2;184;149;95m@[0m[38;2;185;148;95m@[0m[38;2;185;148;94m&[0m[38;2;185;148;93m&[0m[38;2;186;149;96m@[0m[38;2;160;123;75mB[0m[38;2;140;101;57m#[0m[38;2;136;95;56m#[0m[38;2;130;89;54m#[0m[38;2;125;83;50mS[0m[38;2;121;79;47mS[0m[38;2;124;83;50mS[0m[38;2;130;90;55m#[0m[38;2;134;93;59m#[0m[38;2;135;95;62m#[0m[38;2;128;88;54m#[0m[38;2;124;87;54mS[0m[38;2;100;69;39mH[0m[38;2;79;53;32mh[0m[38;2;54;31;20mA[0m[38;2;39;23;12ms[0m");
	$display("[38;2;172;133;78m&[0m[38;2;173;134;79m&[0m[38;2;173;134;78m&[0m[38;2;173;134;79m&[0m[38;2;173;134;78m&[0m[38;2;174;135;78m&[0m[38;2;174;135;78m&[0m[38;2;174;135;76m&[0m[38;2;174;134;76m&[0m[38;2;173;135;77m&[0m[38;2;175;136;79m&[0m[38;2;174;136;79m&[0m[38;2;175;137;79m&[0m[38;2;176;137;80m&[0m[38;2;177;136;80m&[0m[38;2;177;136;80m&[0m[38;2;177;136;80m&[0m[38;2;177;136;80m&[0m[38;2;177;136;80m&[0m[38;2;177;136;81m&[0m[38;2;177;136;81m&[0m[38;2;177;136;81m&[0m[38;2;178;137;82m&[0m[38;2;178;137;80m&[0m[38;2;178;137;80m&[0m[38;2;177;137;79m&[0m[38;2;177;137;79m&[0m[38;2;178;137;79m&[0m[38;2;177;137;79m&[0m[38;2;178;137;79m&[0m[38;2;178;137;79m&[0m[38;2;178;137;79m&[0m[38;2;177;137;79m&[0m[38;2;176;136;78m&[0m[38;2;177;136;78m&[0m[38;2;177;137;78m&[0m[38;2;177;137;78m&[0m[38;2;177;136;78m&[0m[38;2;177;137;78m&[0m[38;2;177;137;78m&[0m[38;2;176;136;77m&[0m[38;2;176;134;78m&[0m[38;2;174;135;78m&[0m[38;2;173;129;82m&[0m[38;2;107;47;29mM[0m[38;2;68;2;3ms[0m[38;2;78;30;16m2[0m[38;2;178;145;120m@[0m[38;2;183;165;131m@[0m[38;2;145;132;93mB[0m[38;2;196;181;143m@[0m[38;2;179;163;128m@[0m[38;2;185;170;132m@[0m[38;2;194;179;140m@[0m[38;2;184;169;130m@[0m[38;2;197;182;145m@[0m[38;2;199;183;153m@[0m[38;2;105;88;61mS[0m[38;2;169;152;120m@[0m[38;2;159;143;110m&[0m[38;2;187;172;134m@[0m[38;2;216;201;165m@[0m[38;2;176;159;127m@[0m[38;2;154;134;103m&[0m[38;2;150;127;97m&[0m[38;2;99;77;50mG[0m[38;2;101;82;54mG[0m[38;2;179;163;128m@[0m[38;2;193;181;140m@[0m[38;2;222;207;171m@[0m[38;2;176;160;128m@[0m[38;2;144;127;97mB[0m[38;2;190;174;141m@[0m[38;2;205;189;154m@[0m[38;2;208;192;158m@[0m[38;2;193;177;141m@[0m[38;2;185;170;132m@[0m[38;2;192;177;138m@[0m[38;2;197;181;141m@[0m[38;2;200;186;146m@[0m[38;2;149;135;103m&[0m[38;2;88;71;50mH[0m[38;2;60;38;26m2[0m[38;2;46;19;12ms[0m[38;2;59;13;11ms[0m[38;2;77;8;11mX[0m[38;2;84;7;9mA[0m[38;2;85;8;6mX[0m[38;2;82;8;5mX[0m[38;2;74;7;5mX[0m[38;2;73;14;7mX[0m[38;2;127;78;49mS[0m[38;2;151;108;62m9[0m[38;2;151;110;61m9[0m[38;2;151;109;61m9[0m[38;2;150;108;60m9[0m[38;2;151;109;61m9[0m[38;2;169;127;79m&[0m[38;2;172;131;83m&[0m[38;2;173;133;84m&[0m[38;2;171;132;83m&[0m[38;2;172;134;86m&[0m[38;2;147;111;67m9[0m[38;2;112;78;39mG[0m[38;2;128;91;53m#[0m[38;2;154;112;70mB[0m[38;2;172;130;82m&[0m[38;2;183;145;92m&[0m[38;2;184;149;93m&[0m[38;2;183;149;93m&[0m[38;2;184;148;95m&[0m[38;2;183;149;94m&[0m[38;2;181;148;94m&[0m[38;2;182;148;94m&[0m[38;2;184;148;94m&[0m[38;2;185;147;95m&[0m[38;2;185;148;95m@[0m[38;2;186;149;96m@[0m[38;2;179;141;93m&[0m[38;2;144;106;63m9[0m[38;2;118;79;44mG[0m[38;2;113;74;42mG[0m[38;2;115;75;45mG[0m[38;2;118;78;49mS[0m[38;2;119;79;50mS[0m[38;2;124;81;52mS[0m[38;2;131;87;57m#[0m[38;2;137;90;61m#[0m[38;2;140;92;63m#[0m[38;2;128;82;53mS[0m[38;2;119;77;46mG[0m[38;2;101;64;35mM[0m[38;2;95;63;40mM[0m[38;2;71;44;27m5[0m[38;2;44;26;14ms[0m");
	$display("[38;2;161;122;72mB[0m[38;2;163;123;73mB[0m[38;2;163;123;74mB[0m[38;2;163;124;74mB[0m[38;2;166;126;76mB[0m[38;2;169;128;78m&[0m[38;2;172;131;80m&[0m[38;2;174;133;80m&[0m[38;2;175;134;78m&[0m[38;2;173;134;78m&[0m[38;2;171;134;78m&[0m[38;2;172;134;79m&[0m[38;2;172;135;79m&[0m[38;2;171;135;79m&[0m[38;2;173;134;80m&[0m[38;2;174;134;79m&[0m[38;2;173;134;79m&[0m[38;2;173;134;79m&[0m[38;2;173;133;78m&[0m[38;2;173;134;78m&[0m[38;2;174;134;78m&[0m[38;2;174;135;79m&[0m[38;2;174;135;79m&[0m[38;2;174;135;80m&[0m[38;2;175;135;80m&[0m[38;2;174;135;80m&[0m[38;2;174;135;80m&[0m[38;2;174;135;80m&[0m[38;2;174;135;80m&[0m[38;2;174;135;79m&[0m[38;2;175;135;80m&[0m[38;2;175;136;80m&[0m[38;2;175;136;80m&[0m[38;2;174;135;79m&[0m[38;2;174;135;79m&[0m[38;2;173;134;78m&[0m[38;2;173;134;78m&[0m[38;2;174;133;78m&[0m[38;2;174;133;79m&[0m[38;2;174;133;79m&[0m[38;2;174;133;78m&[0m[38;2;173;133;78m&[0m[38;2;172;134;76m&[0m[38;2;175;128;82m&[0m[38;2;104;48;30mM[0m[38;2;69;19;11mX[0m[38;2;174;142;114m@[0m[38;2;188;165;132m@[0m[38;2;123;106;73m9[0m[38;2;187;169;135m@[0m[38;2;175;155;120m@[0m[38;2;162;147;110m&[0m[38;2;192;176;139m@[0m[38;2;178;163;124m@[0m[38;2;164;149;110m&[0m[38;2;206;190;153m@[0m[38;2;104;87;58mS[0m[38;2;124;106;81m9[0m[38;2;159;142;111m&[0m[38;2;162;145;109m&[0m[38;2;191;174;135m@[0m[38;2;209;194;161m@[0m[38;2;113;97;70m#[0m[38;2;136;116;86mB[0m[38;2;167;139;104m&[0m[38;2;193;161;122m@[0m[38;2;129;101;72m9[0m[38;2;103;81;59mG[0m[38;2;176;163;127m@[0m[38;2;202;187;149m@[0m[38;2;223;207;173m@[0m[38;2;132;115;84m9[0m[38;2;146;130;99m&[0m[38;2;190;175;140m@[0m[38;2;205;190;149m@[0m[38;2;197;182;142m@[0m[38;2;186;171;133m@[0m[38;2;177;161;125m@[0m[38;2;190;174;137m@[0m[38;2;192;176;134m@[0m[38;2;205;186;144m@[0m[38;2;161;142;108m&[0m[38;2;121;102;77m9[0m[38;2;102;87;64mS[0m[38;2;58;41;24m2[0m[38;2;46;16;9mr[0m[38;2;66;10;12mX[0m[38;2;80;7;8mX[0m[38;2;78;7;6mX[0m[38;2;76;5;9mX[0m[38;2;70;3;8ms[0m[38;2;83;25;16m2[0m[38;2;140;96;56m#[0m[38;2;148;108;58m9[0m[38;2;147;107;58m9[0m[38;2;146;106;57m9[0m[38;2;147;107;58m9[0m[38;2;165;125;76mB[0m[38;2;171;131;82m&[0m[38;2;171;132;83m&[0m[38;2;170;132;83m&[0m[38;2;171;133;85m&[0m[38;2;146;112;67m9[0m[38;2;110;78;40mG[0m[38;2;126;90;52mS[0m[38;2;151;110;68m9[0m[38;2;170;127;82m&[0m[38;2;182;142;93m&[0m[38;2;183;147;94m&[0m[38;2;183;146;95m&[0m[38;2;183;146;95m&[0m[38;2;183;147;94m&[0m[38;2;183;147;93m&[0m[38;2;183;147;93m&[0m[38;2;184;145;93m&[0m[38;2;186;146;95m&[0m[38;2;182;142;93m&[0m[38;2;163;122;79mB[0m[38;2;144;102;65m9[0m[38;2;134;91;57m#[0m[38;2;129;85;54mS[0m[38;2;130;86;54m#[0m[38;2;124;80;48mS[0m[38;2;125;80;50mS[0m[38;2;125;81;51mS[0m[38;2;126;81;52mS[0m[38;2;131;87;58m#[0m[38;2;136;93;61m#[0m[38;2;139;97;61m#[0m[38;2;146;103;67m9[0m[38;2;162;119;78mB[0m[38;2;178;136;89m&[0m[38;2;182;141;93m&[0m[38;2;172;131;87m&[0m[38;2;138;100;65m9[0m");
	$display("[38;2;106;76;49mG[0m[38;2;110;78;53mG[0m[38;2;112;78;52mG[0m[38;2;114;81;51mS[0m[38;2;115;83;52mS[0m[38;2;116;82;54mS[0m[38;2;120;86;56mS[0m[38;2;129;93;59m#[0m[38;2;137;101;62m9[0m[38;2;150;114;70mB[0m[38;2;163;125;76mB[0m[38;2;169;131;75m&[0m[38;2;169;132;75m&[0m[38;2;168;132;77m&[0m[38;2;169;131;81m&[0m[38;2;171;132;78m&[0m[38;2;171;132;76m&[0m[38;2;172;131;77m&[0m[38;2;172;132;77m&[0m[38;2;172;133;78m&[0m[38;2;172;133;78m&[0m[38;2;172;133;77m&[0m[38;2;172;133;77m&[0m[38;2;172;133;78m&[0m[38;2;173;134;79m&[0m[38;2;173;134;79m&[0m[38;2;172;133;78m&[0m[38;2;172;133;78m&[0m[38;2;172;133;78m&[0m[38;2;173;134;79m&[0m[38;2;172;133;78m&[0m[38;2;172;133;78m&[0m[38;2;172;133;78m&[0m[38;2;173;134;79m&[0m[38;2;173;134;79m&[0m[38;2;172;133;78m&[0m[38;2;171;132;77m&[0m[38;2;172;131;77m&[0m[38;2;172;131;77m&[0m[38;2;172;131;77m&[0m[38;2;172;131;77m&[0m[38;2;170;130;78m&[0m[38;2;170;130;71mB[0m[38;2;173;129;75m&[0m[38;2;125;83;53mS[0m[38;2;144;111;84mB[0m[38;2;193;173;141m@[0m[38;2;106;89;59mS[0m[38;2;155;140;110m&[0m[38;2;172;155;124m@[0m[38;2;123;105;72m9[0m[38;2;175;158;120m@[0m[38;2;185;168;132m@[0m[38;2;137;120;86mB[0m[38;2;178;160;128m@[0m[38;2;132;114;84m9[0m[38;2;70;51;25m5[0m[38;2;163;145;119m&[0m[38;2;126;109;77m9[0m[38;2;178;162;123m@[0m[38;2;188;173;132m@[0m[38;2;182;165;131m@[0m[38;2;74;59;34mh[0m[38;2;129;111;83m9[0m[38;2;161;132;96m&[0m[38;2;196;161;120m@[0m[38;2;202;172;130m@[0m[38;2;132;108;73m9[0m[38;2;104;87;61mS[0m[38;2;179;164;131m@[0m[38;2;212;197;156m@[0m[38;2;193;177;142m@[0m[38;2;96;79;50mG[0m[38;2;168;152;118m@[0m[38;2;189;174;133m@[0m[38;2;191;176;136m@[0m[38;2;190;175;137m@[0m[38;2;161;145;110m&[0m[38;2;177;162;127m@[0m[38;2;179;164;128m@[0m[38;2;187;171;132m@[0m[38;2;200;184;149m@[0m[38;2;133;117;87mB[0m[38;2;129;111;82m9[0m[38;2;156;142;108m&[0m[38;2;106;93;68mS[0m[38;2;56;29;19mA[0m[38;2;54;9;4mr[0m[38;2;66;8;7ms[0m[38;2;72;5;7ms[0m[38;2;76;5;6mX[0m[38;2;73;7;2ms[0m[38;2;114;65;37mH[0m[38;2;147;106;60m9[0m[38;2;146;105;56m9[0m[38;2;146;104;58m9[0m[38;2;146;105;56m9[0m[38;2;162;124;74mB[0m[38;2;169;131;82m&[0m[38;2;169;131;82m&[0m[38;2;169;131;82m&[0m[38;2;170;132;83m&[0m[38;2;144;109;66m9[0m[38;2;106;76;42mG[0m[38;2;125;87;54mS[0m[38;2;152;110;68m9[0m[38;2;170;126;82m&[0m[38;2;181;139;93m&[0m[38;2;182;144;95m&[0m[38;2;183;145;96m&[0m[38;2;183;144;96m&[0m[38;2;182;144;95m&[0m[38;2;182;145;92m&[0m[38;2;183;146;92m&[0m[38;2;182;145;94m&[0m[38;2;171;132;88m&[0m[38;2;147;105;66m9[0m[38;2;139;97;58m#[0m[38;2;147;104;68m9[0m[38;2;150;106;71m9[0m[38;2;148;102;66m9[0m[38;2;148;102;69m9[0m[38;2;144;99;67m9[0m[38;2;142;97;65m9[0m[38;2;139;95;63m#[0m[38;2;144;99;66m9[0m[38;2;159;115;78mB[0m[38;2;172;131;89m&[0m[38;2;182;142;95m&[0m[38;2;185;145;96m&[0m[38;2;185;144;96m&[0m[38;2;184;143;94m&[0m[38;2;183;143;94m&[0m[38;2;183;142;93m&[0m[38;2;177;136;87m&[0m");
	$display("[38;2;105;75;49mG[0m[38;2;111;77;53mG[0m[38;2;119;83;60mS[0m[38;2;122;87;60mS[0m[38;2;121;87;59mS[0m[38;2;117;84;58mS[0m[38;2;114;81;56mS[0m[38;2;111;78;53mG[0m[38;2;108;76;47mG[0m[38;2;111;77;48mG[0m[38;2;125;90;55m#[0m[38;2;142;104;62m9[0m[38;2;158;121;74mB[0m[38;2;166;129;81m&[0m[38;2;167;130;78m&[0m[38;2;169;129;75m&[0m[38;2;169;130;74m&[0m[38;2;170;129;75m&[0m[38;2;169;129;77m&[0m[38;2;169;129;77m&[0m[38;2;169;129;77m&[0m[38;2;169;129;78m&[0m[38;2;169;129;78m&[0m[38;2;169;130;77m&[0m[38;2;170;130;77m&[0m[38;2;170;130;77m&[0m[38;2;170;130;77m&[0m[38;2;170;130;77m&[0m[38;2;170;130;77m&[0m[38;2;171;131;78m&[0m[38;2;170;131;78m&[0m[38;2;169;130;77m&[0m[38;2;169;130;77m&[0m[38;2;169;130;77m&[0m[38;2;169;129;76m&[0m[38;2;169;129;76m&[0m[38;2;168;129;76m&[0m[38;2;170;129;76m&[0m[38;2;170;129;76m&[0m[38;2;170;129;76m&[0m[38;2;170;129;76m&[0m[38;2;170;128;75m&[0m[38;2;168;127;74mB[0m[38;2;164;127;77mB[0m[38;2;155;127;83mB[0m[38;2;183;164;125m@[0m[38;2;125;109;83m9[0m[38;2;100;84;59mG[0m[38;2;171;153;128m@[0m[38;2;107;89;65mS[0m[38;2;108;92;64mS[0m[38;2;183;168;130m@[0m[38;2;155;138;105m&[0m[38;2;117;99;71m#[0m[38;2;154;136;111m&[0m[38;2;54;36;16mA[0m[38;2;108;91;70mS[0m[38;2;132;116;90mB[0m[38;2;124;108;75m9[0m[38;2;183;169;132m@[0m[38;2;182;168;129m@[0m[38;2;150;131;99m&[0m[38;2;82;63;39mM[0m[38;2;136;118;89mB[0m[38;2;156;130;94m&[0m[38;2;194;160;121m@[0m[38;2;204;170;123m@[0m[38;2;201;171;127m@[0m[38;2;127;105;73m9[0m[38;2;111;93;66m#[0m[38;2;184;169;131m@[0m[38;2;210;195;156m@[0m[38;2;123;106;78m9[0m[38;2;103;86;59mS[0m[38;2;184;168;133m@[0m[38;2;186;170;131m@[0m[38;2;186;172;132m@[0m[38;2;174;158;123m@[0m[38;2;145;129;97mB[0m[38;2;172;155;124m@[0m[38;2;148;132;98m&[0m[38;2;188;172;135m@[0m[38;2;192;177;139m@[0m[38;2;102;84;56mG[0m[38;2;136;113;84mB[0m[38;2;184;166;126m@[0m[38;2;158;145;109m&[0m[38;2;83;64;43mM[0m[38;2;52;15;8ms[0m[38;2;65;8;7ms[0m[38;2;76;6;8mX[0m[38;2;76;5;5mX[0m[38;2;91;40;22m3[0m[38;2;141;100;61m9[0m[38;2;142;103;53m#[0m[38;2;143;103;56m9[0m[38;2;143;104;55m9[0m[38;2;160;122;73mB[0m[38;2;168;130;81m&[0m[38;2;168;130;81m&[0m[38;2;168;130;81m&[0m[38;2;169;130;81m&[0m[38;2;143;108;65m9[0m[38;2;105;75;41mH[0m[38;2;124;86;53mS[0m[38;2;150;108;66m9[0m[38;2;167;124;79mB[0m[38;2;178;139;92m&[0m[38;2;180;144;95m&[0m[38;2;181;145;95m&[0m[38;2;180;143;93m&[0m[38;2;180;142;91m&[0m[38;2;180;143;90m&[0m[38;2;180;143;93m&[0m[38;2;161;123;80mB[0m[38;2;140;99;62m9[0m[38;2;146;102;68m9[0m[38;2;158;114;77mB[0m[38;2;164;119;81mB[0m[38;2;158;113;74mB[0m[38;2;149;104;66m9[0m[38;2;149;104;68m9[0m[38;2;147;103;69m9[0m[38;2;148;104;68m9[0m[38;2;157;114;76mB[0m[38;2;174;130;92m&[0m[38;2;185;142;101m@[0m[38;2;186;145;99m@[0m[38;2;186;145;96m&[0m[38;2;184;146;95m&[0m[38;2;182;143;94m&[0m[38;2;182;143;94m&[0m[38;2;181;142;93m&[0m[38;2;179;140;92m&[0m[38;2;172;131;85m&[0m");
	$display("[38;2;158;117;86mB[0m[38;2;144;104;74m9[0m[38;2;129;92;64m#[0m[38;2;119;83;57mS[0m[38;2;116;83;57mS[0m[38;2;117;85;58mS[0m[38;2;119;85;58mS[0m[38;2;125;91;61m#[0m[38;2;126;91;58m#[0m[38;2;125;90;56m#[0m[38;2;122;86;57mS[0m[38;2;121;84;57mS[0m[38;2;125;88;56mS[0m[38;2;140;104;64m9[0m[38;2;160;124;75mB[0m[38;2;168;129;73mB[0m[38;2;168;127;74mB[0m[38;2;168;127;76mB[0m[38;2;167;127;75mB[0m[38;2;168;126;76mB[0m[38;2;167;126;76mB[0m[38;2;167;126;76mB[0m[38;2;167;126;76mB[0m[38;2;166;127;75mB[0m[38;2;166;127;75mB[0m[38;2;166;127;75mB[0m[38;2;167;128;76mB[0m[38;2;168;128;76m&[0m[38;2;168;128;76m&[0m[38;2;168;128;76m&[0m[38;2;168;128;75mB[0m[38;2;167;128;74mB[0m[38;2;167;127;75mB[0m[38;2;167;127;75mB[0m[38;2;167;126;75mB[0m[38;2;167;127;75mB[0m[38;2;168;127;75mB[0m[38;2;168;127;75mB[0m[38;2;167;126;74mB[0m[38;2;167;126;74mB[0m[38;2;167;126;74mB[0m[38;2;168;125;74mB[0m[38;2;168;126;76mB[0m[38;2;155;122;77mB[0m[38;2;169;145;105m&[0m[38;2;166;146;115m&[0m[38;2;71;54;33m3[0m[38;2;132;116;91mB[0m[38;2;117;100;80m#[0m[38;2;50;35;16mA[0m[38;2;137;124;95mB[0m[38;2;178;163;129m@[0m[38;2;103;89;61mS[0m[38;2;129;117;88mB[0m[38;2;75;61;42mh[0m[38;2;53;37;22mA[0m[38;2;127;112;88m9[0m[38;2;73;58;33mh[0m[38;2;140;125;99mB[0m[38;2;181;166;129m@[0m[38;2;176;161;123m@[0m[38;2;114;91;64mS[0m[38;2;121;96;71m#[0m[38;2;148;124;93mB[0m[38;2;149;123;89mB[0m[38;2;195;163;124m@[0m[38;2;203;168;123m@[0m[38;2;202;170;126m@[0m[38;2;194;169;125m@[0m[38;2;120;99;62m#[0m[38;2;120;100;72m#[0m[38;2;190;174;139m@[0m[38;2;167;151;117m@[0m[38;2;70;52;33m3[0m[38;2;152;136;107m&[0m[38;2;185;169;132m@[0m[38;2;183;168;127m@[0m[38;2;186;170;134m@[0m[38;2;132;115;84m9[0m[38;2;170;154;123m@[0m[38;2;131;114;83m9[0m[38;2;149;133;99m&[0m[38;2;192;177;136m@[0m[38;2;164;148;116m@[0m[38;2;79;60;38mh[0m[38;2;146;132;98m&[0m[38;2;186;173;129m@[0m[38;2;181;166;128m@[0m[38;2;104;84;60mS[0m[38;2;59;18;13mX[0m[38;2;73;8;9mX[0m[38;2;74;6;8mX[0m[38;2;78;28;18m2[0m[38;2;136;94;59m#[0m[38;2;140;101;53m#[0m[38;2;140;102;54m#[0m[38;2;140;102;54m#[0m[38;2;159;121;73mB[0m[38;2;167;129;81m&[0m[38;2;166;128;80m&[0m[38;2;167;129;81m&[0m[38;2;167;129;81m&[0m[38;2;141;109;63m9[0m[38;2;102;74;39mH[0m[38;2;120;84;50mS[0m[38;2;146;107;65m9[0m[38;2;165;124;78mB[0m[38;2;176;138;91m&[0m[38;2;179;143;94m&[0m[38;2;179;143;93m&[0m[38;2;179;143;92m&[0m[38;2;180;144;92m&[0m[38;2;177;140;92m&[0m[38;2;153;114;71mB[0m[38;2;138;99;59m#[0m[38;2;152;110;71mB[0m[38;2;162;118;79mB[0m[38;2;164;119;80mB[0m[38;2;164;119;80mB[0m[38;2;156;112;72mB[0m[38;2;148;102;63m9[0m[38;2;147;102;64m9[0m[38;2;154;110;70mB[0m[38;2;169;126;85m&[0m[38;2;182;139;97m&[0m[38;2;184;141;98m&[0m[38;2;183;141;96m&[0m[38;2;182;142;97m&[0m[38;2;183;143;99m&[0m[38;2;183;143;100m&[0m[38;2;183;142;98m&[0m[38;2;182;142;96m&[0m[38;2;182;141;95m&[0m[38;2;180;139;93m&[0m[38;2;181;140;93m&[0m");
	$display("[38;2;167;125;94m&[0m[38;2;169;128;95m&[0m[38;2;167;129;95m&[0m[38;2;158;121;90mB[0m[38;2;138;103;74m9[0m[38;2;124;90;60m#[0m[38;2;129;93;62m#[0m[38;2;145;106;74m9[0m[38;2;148;106;73m9[0m[38;2;147;106;70m9[0m[38;2;141;101;67m9[0m[38;2;131;93;62m#[0m[38;2;122;86;56mS[0m[38;2;120;85;52mS[0m[38;2;127;91;56m#[0m[38;2;151;113;71mB[0m[38;2;163;125;77mB[0m[38;2;163;125;73mB[0m[38;2;165;124;74mB[0m[38;2;165;124;76mB[0m[38;2;165;124;75mB[0m[38;2;164;125;74mB[0m[38;2;164;125;74mB[0m[38;2;165;125;74mB[0m[38;2;165;125;74mB[0m[38;2;166;125;75mB[0m[38;2;166;126;77mB[0m[38;2;167;126;77mB[0m[38;2;166;126;74mB[0m[38;2;166;125;74mB[0m[38;2;165;125;74mB[0m[38;2;165;125;72mB[0m[38;2;165;125;72mB[0m[38;2;165;125;72mB[0m[38;2;165;125;72mB[0m[38;2;165;125;72mB[0m[38;2;164;125;72mB[0m[38;2;164;125;72mB[0m[38;2;164;124;71mB[0m[38;2;164;124;71mB[0m[38;2;164;124;71mB[0m[38;2;164;124;72mB[0m[38;2;161;124;74mB[0m[38;2;151;125;79mB[0m[38;2;177;159;123m@[0m[38;2;114;99;73m#[0m[38;2;62;52;35m3[0m[38;2;105;94;74m#[0m[38;2;50;35;23mA[0m[38;2;60;43;28m5[0m[38;2;161;144;112m&[0m[38;2;151;132;104m&[0m[38;2;85;68;51mH[0m[38;2;97;82;61mG[0m[38;2;45;28;17mX[0m[38;2;79;62;52mM[0m[38;2;82;67;50mM[0m[38;2;56;41;23m2[0m[38;2;134;118;91mB[0m[38;2;183;166;130m@[0m[38;2;149;134;100m&[0m[38;2;100;79;53mG[0m[38;2;156;130;101m&[0m[38;2;142;118;88mB[0m[38;2;141;117;86mB[0m[38;2;194;164;124m@[0m[38;2;199;167;121m@[0m[38;2;202;168;124m@[0m[38;2;203;170;121m@[0m[38;2;196;167;119m@[0m[38;2;116;90;58mS[0m[38;2;131;112;80m9[0m[38;2;179;164;130m@[0m[38;2;88;72;50mH[0m[38;2;103;88;62mS[0m[38;2;182;166;132m@[0m[38;2;181;167;127m@[0m[38;2;185;169;133m@[0m[38;2;142;125;92mB[0m[38;2;144;128;93mB[0m[38;2;168;152;120m@[0m[38;2;98;81;52mG[0m[38;2;170;154;117m@[0m[38;2;191;175;136m@[0m[38;2;104;88;63mS[0m[38;2;93;76;55mG[0m[38;2;173;158;123m@[0m[38;2;189;173;128m@[0m[38;2;175;161;122m@[0m[38;2;93;71;49mH[0m[38;2;64;12;9ms[0m[38;2;72;4;9ms[0m[38;2;84;34;22m5[0m[38;2;135;95;60m#[0m[38;2;136;98;53m#[0m[38;2;137;98;55m#[0m[38;2;137;99;54m#[0m[38;2;156;118;72mB[0m[38;2;166;128;81m&[0m[38;2;165;127;81m&[0m[38;2;166;128;82m&[0m[38;2;166;129;81m&[0m[38;2;141;109;65m9[0m[38;2;100;72;38mH[0m[38;2;117;81;49mS[0m[38;2;143;104;64m9[0m[38;2;162;121;76mB[0m[38;2;175;137;89m&[0m[38;2;177;141;90m&[0m[38;2;178;141;91m&[0m[38;2;178;142;92m&[0m[38;2;174;139;91m&[0m[38;2;146;109;66m9[0m[38;2;140;102;62m9[0m[38;2;154;115;76mB[0m[38;2;160;120;80mB[0m[38;2;161;117;78mB[0m[38;2;162;117;78mB[0m[38;2;163;118;79mB[0m[38;2;156;112;73mB[0m[38;2;151;107;67m9[0m[38;2;169;124;84m&[0m[38;2;180;137;95m&[0m[38;2;182;140;97m&[0m[38;2;182;140;96m&[0m[38;2;181;140;94m&[0m[38;2;180;139;94m&[0m[38;2;181;139;95m&[0m[38;2;181;139;96m&[0m[38;2;181;138;96m&[0m[38;2;182;139;95m&[0m[38;2;181;140;94m&[0m[38;2;182;140;95m&[0m[38;2;178;136;95m&[0m[38;2;163;120;87mB[0m");
	$display("[38;2;165;124;93m&[0m[38;2;168;127;93m&[0m[38;2;170;130;95m&[0m[38;2;170;131;95m&[0m[38;2;170;130;95m&[0m[38;2;165;124;90m&[0m[38;2;157;116;82mB[0m[38;2;148;108;73m9[0m[38;2;146;105;70m9[0m[38;2;147;107;71m9[0m[38;2;147;106;70m9[0m[38;2;146;107;71m9[0m[38;2;141;103;68m9[0m[38;2;131;93;59m#[0m[38;2;121;84;55mS[0m[38;2;118;82;54mS[0m[38;2;135;101;60m#[0m[38;2;159;122;76mB[0m[38;2;173;132;88m&[0m[38;2;178;137;91m&[0m[38;2;177;137;89m&[0m[38;2;175;138;87m&[0m[38;2;174;138;85m&[0m[38;2;173;136;85m&[0m[38;2;171;134;85m&[0m[38;2;167;130;84m&[0m[38;2;150;113;70mB[0m[38;2;150;112;67m9[0m[38;2;161;122;73mB[0m[38;2;162;123;73mB[0m[38;2;163;124;73mB[0m[38;2;162;123;72mB[0m[38;2;162;123;73mB[0m[38;2;161;122;73mB[0m[38;2;160;122;72mB[0m[38;2;161;122;72mB[0m[38;2;161;123;73mB[0m[38;2;161;122;73mB[0m[38;2;160;121;71mB[0m[38;2;160;121;72mB[0m[38;2;160;121;72mB[0m[38;2;160;121;72mB[0m[38;2;155;120;72mB[0m[38;2;157;133;90m&[0m[38;2;168;151;120m@[0m[38;2;68;54;35m3[0m[38;2;55;41;31m2[0m[38;2;47;34;21mA[0m[38;2;54;35;26m2[0m[38;2;107;87;70mS[0m[38;2;159;143;110m&[0m[38;2;89;72;55mH[0m[38;2;68;51;43m3[0m[38;2;50;35;22mA[0m[38;2;48;33;22mA[0m[38;2;65;50;40m3[0m[38;2;44;31;22mX[0m[38;2;50;36;22mA[0m[38;2;141;125;94mB[0m[38;2;178;160;127m@[0m[38;2;98;80;53mG[0m[38;2;131;106;77m9[0m[38;2;167;139;109m&[0m[38;2;130;102;76m9[0m[38;2;134;106;79m9[0m[38;2;179;151;113m@[0m[38;2;174;146;106m&[0m[38;2;173;142;104m&[0m[38;2;176;145;104m&[0m[38;2;181;150;107m@[0m[38;2;175;147;112m@[0m[38;2;99;76;49mG[0m[38;2;148;130;103m&[0m[38;2;121;104;78m9[0m[38;2;68;52;31m3[0m[38;2;169;153;121m@[0m[38;2;182;166;127m@[0m[38;2;183;166;129m@[0m[38;2;151;133;105m&[0m[38;2;106;89;63mS[0m[38;2;182;165;132m@[0m[38;2;117;99;74m#[0m[38;2;108;92;64mS[0m[38;2;182;167;130m@[0m[38;2;152;137;103m&[0m[38;2;64;48;27m5[0m[38;2;144;128;104m&[0m[38;2;184;167;128m@[0m[38;2;187;172;129m@[0m[38;2;166;145;112m&[0m[38;2;75;32;25m5[0m[38;2;57;4;3mr[0m[38;2;103;62;37mH[0m[38;2;134;98;57m#[0m[38;2;134;97;53m#[0m[38;2;135;97;54m#[0m[38;2;137;98;54m#[0m[38;2;155;116;72mB[0m[38;2;165;127;82m&[0m[38;2;165;126;81m&[0m[38;2;165;126;82m&[0m[38;2;166;128;81m&[0m[38;2;141;109;66m9[0m[38;2;99;72;39mH[0m[38;2;115;79;49mG[0m[38;2;141;101;63m9[0m[38;2;159;118;76mB[0m[38;2;173;135;85m&[0m[38;2;175;140;85m&[0m[38;2;177;142;92m&[0m[38;2;171;134;88m&[0m[38;2;144;104;62m9[0m[38;2;144;103;65m9[0m[38;2;160;117;82mB[0m[38;2;162;119;83mB[0m[38;2;160;117;79mB[0m[38;2;160;117;78mB[0m[38;2;160;115;77mB[0m[38;2;161;117;78mB[0m[38;2;168;124;85m&[0m[38;2;178;136;94m&[0m[38;2;182;140;97m&[0m[38;2;180;139;95m&[0m[38;2;180;139;94m&[0m[38;2;179;139;95m&[0m[38;2;178;139;95m&[0m[38;2;179;138;95m&[0m[38;2;179;139;93m&[0m[38;2;180;139;90m&[0m[38;2;181;137;90m&[0m[38;2;181;138;92m&[0m[38;2;176;135;93m&[0m[38;2;157;117;84mB[0m[38;2;122;83;57mS[0m[38;2;105;68;45mH[0m");
	$display("[38;2;163;123;88m&[0m[38;2;164;124;89m&[0m[38;2;166;125;90m&[0m[38;2;166;126;91m&[0m[38;2;166;126;91m&[0m[38;2;168;128;92m&[0m[38;2;168;128;93m&[0m[38;2;165;125;90m&[0m[38;2;157;117;82mB[0m[38;2;147;107;72m9[0m[38;2;144;104;69m9[0m[38;2;145;105;70m9[0m[38;2;145;105;70m9[0m[38;2;145;105;70m9[0m[38;2;139;100;65m9[0m[38;2;127;91;59m#[0m[38;2;117;82;50mS[0m[38;2;129;91;56m#[0m[38;2;173;132;93m&[0m[38;2;191;152;102m@[0m[38;2;186;148;96m@[0m[38;2;183;145;97m&[0m[38;2;181;144;95m&[0m[38;2;180;143;94m&[0m[38;2;168;131;86m&[0m[38;2;149;113;74mB[0m[38;2;135;101;64m9[0m[38;2;119;84;45mS[0m[38;2;151;113;68mB[0m[38;2;157;119;71mB[0m[38;2;157;120;69mB[0m[38;2;158;120;71mB[0m[38;2;157;120;71mB[0m[38;2;157;119;70mB[0m[38;2;158;120;71mB[0m[38;2;158;120;71mB[0m[38;2;157;119;70mB[0m[38;2;157;119;69mB[0m[38;2;157;119;69mB[0m[38;2;157;119;69mB[0m[38;2;157;119;69mB[0m[38;2;157;120;69mB[0m[38;2;149;116;67mB[0m[38;2;165;141;98m&[0m[38;2;143;126;98mB[0m[38;2;45;30;18mX[0m[38;2;40;26;19ms[0m[38;2;42;28;16mX[0m[38;2;98;75;59mG[0m[38;2;134;113;89mB[0m[38;2;123;112;86m9[0m[38;2;45;31;18mX[0m[38;2;45;28;22mX[0m[38;2;46;29;21mX[0m[38;2;45;29;21mX[0m[38;2;45;29;23mX[0m[38;2;41;28;20mX[0m[38;2;65;52;32m3[0m[38;2;169;149;121m@[0m[38;2;127;106;83m9[0m[38;2;76;54;34mh[0m[38;2;183;152;110m@[0m[38;2;168;141;103m&[0m[38;2;108;83;59mS[0m[38;2;153;121;90mB[0m[38;2;199;166;124m@[0m[38;2;196;164;119m@[0m[38;2;193;161;116m@[0m[38;2;190;158;114m@[0m[38;2;185;153;107m@[0m[38;2;178;148;106m@[0m[38;2;152;124;90mB[0m[38;2;96;75;50mH[0m[38;2;122;106;88m9[0m[38;2;54;38;24m2[0m[38;2;143;126;98mB[0m[38;2;182;164;126m@[0m[38;2;181;164;125m@[0m[38;2;154;138;105m&[0m[38;2;58;42;27m2[0m[38;2;134;117;90mB[0m[38;2;165;145;115m&[0m[38;2;69;54;35m3[0m[38;2;145;132;101m&[0m[38;2;172;156;123m@[0m[38;2;73;59;38mh[0m[38;2;98;84;62mG[0m[38;2;178;162;124m@[0m[38;2;184;170;123m@[0m[38;2;183;167;126m@[0m[38;2;130;103;79m9[0m[38;2;78;40;23m5[0m[38;2;128;92;56m#[0m[38;2;131;98;54m#[0m[38;2;131;97;52m#[0m[38;2;133;96;52m#[0m[38;2;134;95;53m#[0m[38;2;153;113;70mB[0m[38;2;163;124;80mB[0m[38;2;163;124;80mB[0m[38;2;163;124;79mB[0m[38;2;163;125;78mB[0m[38;2;140;109;67m9[0m[38;2;97;71;38mH[0m[38;2;111;77;46mG[0m[38;2;139;100;61m9[0m[38;2;156;117;74mB[0m[38;2;169;133;81m&[0m[38;2;173;137;87m&[0m[38;2;166;128;88m&[0m[38;2;137;100;62m9[0m[38;2;144;103;68m9[0m[38;2;159;115;80mB[0m[38;2;160;116;79mB[0m[38;2;160;116;78mB[0m[38;2;159;116;79mB[0m[38;2;159;115;79mB[0m[38;2;165;121;83mB[0m[38;2;176;132;92m&[0m[38;2;182;138;97m&[0m[38;2;180;138;95m&[0m[38;2;180;138;96m&[0m[38;2;179;138;95m&[0m[38;2;179;138;94m&[0m[38;2;179;138;94m&[0m[38;2;179;138;94m&[0m[38;2;178;139;91m&[0m[38;2;179;139;91m&[0m[38;2;181;138;91m&[0m[38;2;172;130;88m&[0m[38;2;147;108;72m9[0m[38;2;114;78;50mG[0m[38;2;101;65;42mH[0m[38;2;110;73;49mG[0m[38;2;125;84;54mS[0m");
	$display("[38;2;161;121;86mB[0m[38;2;162;121;86mB[0m[38;2;163;123;88m&[0m[38;2;163;123;88m&[0m[38;2;164;124;89m&[0m[38;2;165;125;90m&[0m[38;2;165;125;90m&[0m[38;2;166;126;91m&[0m[38;2;167;127;92m&[0m[38;2;164;124;89m&[0m[38;2;154;114;79mB[0m[38;2;144;104;69m9[0m[38;2;142;102;67m9[0m[38;2;144;103;68m9[0m[38;2;145;103;68m9[0m[38;2;143;103;70m9[0m[38;2;135;96;65m#[0m[38;2;121;82;54mS[0m[38;2;131;93;63m#[0m[38;2;169;132;91m&[0m[38;2;183;147;96m&[0m[38;2;185;147;98m@[0m[38;2;183;145;95m&[0m[38;2;183;145;96m&[0m[38;2;164;127;82m&[0m[38;2;141;107;67m9[0m[38;2;131;100;62m#[0m[38;2;113;81;41mG[0m[38;2;148;109;64m9[0m[38;2;156;118;70mB[0m[38;2;156;118;67mB[0m[38;2;155;117;68mB[0m[38;2;155;117;68mB[0m[38;2;155;117;68mB[0m[38;2;155;117;68mB[0m[38;2;155;117;68mB[0m[38;2;154;116;67mB[0m[38;2;154;116;68mB[0m[38;2;154;116;68mB[0m[38;2;154;116;68mB[0m[38;2;154;116;68mB[0m[38;2;154;117;70mB[0m[38;2;146;114;70m9[0m[38;2;170;149;110m@[0m[38;2;114;101;76m#[0m[38;2;34;25;15ms[0m[38;2;38;24;17ms[0m[38;2;101;73;55mG[0m[38;2;160;131;99m&[0m[38;2;141;120;92mB[0m[38;2;74;57;39mh[0m[38;2;39;24;13ms[0m[38;2;46;26;21mX[0m[38;2;63;40;31m5[0m[38;2;82;59;48mM[0m[38;2;63;42;31m5[0m[38;2;46;32;18mX[0m[38;2;94;79;60mG[0m[38;2;134;112;91mB[0m[38;2;56;34;20mA[0m[38;2;125;101;79m9[0m[38;2;199;165;124m@[0m[38;2;160;129;96m&[0m[38;2;97;68;47mH[0m[38;2;173;139;108m&[0m[38;2;198;164;120m@[0m[38;2;197;164;118m@[0m[38;2;197;164;117m@[0m[38;2;198;164;119m@[0m[38;2;198;165;118m@[0m[38;2;199;165;116m@[0m[38;2;200;165;122m@[0m[38;2;152;123;93mB[0m[38;2;85;64;47mM[0m[38;2;50;36;23mA[0m[38;2;113;97;73m#[0m[38;2;177;161;127m@[0m[38;2;178;163;123m@[0m[38;2;154;139;104m&[0m[38;2;88;76;52mH[0m[38;2;59;46;33m5[0m[38;2;151;136;107m&[0m[38;2;102;89;65mS[0m[38;2;82;69;46mM[0m[38;2;174;156;126m@[0m[38;2;97;81;57mG[0m[38;2;68;53;32m3[0m[38;2;168;153;119m@[0m[38;2;178;165;119m@[0m[38;2;178;166;121m@[0m[38;2;172;153;115m@[0m[38;2;129;102;64m#[0m[38;2;128;97;52m#[0m[38;2;129;97;51m#[0m[38;2;129;95;53m#[0m[38;2;129;94;52m#[0m[38;2;130;93;50m#[0m[38;2;148;111;67m9[0m[38;2;160;122;77mB[0m[38;2;161;123;78mB[0m[38;2;161;124;78mB[0m[38;2;161;124;77mB[0m[38;2;139;107;66m9[0m[38;2;95;69;38mH[0m[38;2;110;75;47mG[0m[38;2;138;98;61m#[0m[38;2;152;115;74mB[0m[38;2;167;131;86m&[0m[38;2;158;121;80mB[0m[38;2;133;93;60m#[0m[38;2;141;102;67m9[0m[38;2;157;116;80mB[0m[38;2;159;115;80mB[0m[38;2;158;114;77mB[0m[38;2;157;114;76mB[0m[38;2;160;117;80mB[0m[38;2;171;128;89m&[0m[38;2;179;137;97m&[0m[38;2;180;138;96m&[0m[38;2;179;138;94m&[0m[38;2;179;138;94m&[0m[38;2;179;138;95m&[0m[38;2;179;137;95m&[0m[38;2;178;136;94m&[0m[38;2;180;138;94m&[0m[38;2;180;138;94m&[0m[38;2;177;134;93m&[0m[38;2;160;119;84mB[0m[38;2;133;94;65m#[0m[38;2;106;68;44mH[0m[38;2;99;60;38mM[0m[38;2;112;73;50mG[0m[38;2;125;83;55mS[0m[38;2;129;85;52mS[0m[38;2;135;90;55m#[0m");
	$display("[38;2;145;108;80mB[0m[38;2;158;118;87mB[0m[38;2;162;119;86mB[0m[38;2;163;119;85mB[0m[38;2;163;120;86mB[0m[38;2;163;122;88m&[0m[38;2;163;122;90m&[0m[38;2;163;123;89m&[0m[38;2;163;125;88m&[0m[38;2;164;124;89m&[0m[38;2;166;126;91m&[0m[38;2;161;121;86mB[0m[38;2;152;112;77mB[0m[38;2;144;103;69m9[0m[38;2;144;100;67m9[0m[38;2;145;102;70m9[0m[38;2;143;103;72m9[0m[38;2;136;99;69m9[0m[38;2;127;89;63m#[0m[38;2;128;91;60m#[0m[38;2;162;128;84m&[0m[38;2;186;150;99m@[0m[38;2;185;148;95m@[0m[38;2;185;148;96m@[0m[38;2;161;125;80mB[0m[38;2;138;104;65m9[0m[38;2;128;97;58m#[0m[38;2;111;79;40mG[0m[38;2;146;109;64m9[0m[38;2;152;116;65mB[0m[38;2;153;116;68mB[0m[38;2;153;115;66mB[0m[38;2;153;115;66mB[0m[38;2;154;115;66mB[0m[38;2;154;115;67mB[0m[38;2;153;114;66mB[0m[38;2;152;114;66mB[0m[38;2;151;113;68mB[0m[38;2;151;113;68mB[0m[38;2;151;113;68mB[0m[38;2;151;113;68mB[0m[38;2;151;113;67m9[0m[38;2;145;110;74m9[0m[38;2;171;149;114m@[0m[38;2;88;79;55mG[0m[38;2;33;20;14mr[0m[38;2;80;53;41mh[0m[38;2;180;145;107m@[0m[38;2;179;145;101m&[0m[38;2;144;114;89mB[0m[38;2;72;47;31m3[0m[38;2;75;52;38mh[0m[38;2;98;71;50mH[0m[38;2;166;134;106m&[0m[38;2;138;102;74m9[0m[38;2;167;133;101m&[0m[38;2;155;124;90mB[0m[38;2;153;121;89mB[0m[38;2;136;104;74m9[0m[38;2;129;97;68m#[0m[38;2;186;156;114m@[0m[38;2;196;163;122m@[0m[38;2;167;133;99m&[0m[38;2;142;108;75m9[0m[38;2;189;155;117m@[0m[38;2;194;161;119m@[0m[38;2;195;163;119m@[0m[38;2;195;163;119m@[0m[38;2;195;163;119m@[0m[38;2;196;162;118m@[0m[38;2;197;163;118m@[0m[38;2;197;162;116m@[0m[38;2;195;163;122m@[0m[38;2;117;95;66m#[0m[38;2;41;25;10ms[0m[38;2;92;77;60mG[0m[38;2;175;158;121m@[0m[38;2;178;162;121m@[0m[38;2;145;131;101m&[0m[38;2;102;90;67mS[0m[38;2;68;56;43mh[0m[38;2;66;54;35m3[0m[38;2;128;118;93mB[0m[38;2;54;42;25m2[0m[38;2;139;120;98mB[0m[38;2;114;97;73m#[0m[38;2;50;35;21mA[0m[38;2;151;137;107m&[0m[38;2;177;161;122m@[0m[38;2;177;161;120m@[0m[38;2;180;160;120m@[0m[38;2;146;121;84mB[0m[38;2;124;94;52m#[0m[38;2;127;94;51m#[0m[38;2;125;92;51mS[0m[38;2;126;91;51mS[0m[38;2;128;90;51mS[0m[38;2;146;109;67m9[0m[38;2;159;122;78mB[0m[38;2;160;123;78mB[0m[38;2;161;124;79mB[0m[38;2;162;124;79mB[0m[38;2;140;108;65m9[0m[38;2;93;69;34mM[0m[38;2;108;75;45mG[0m[38;2;135;97;61m#[0m[38;2;150;112;75mB[0m[38;2;147;108;71m9[0m[38;2;131;92;56m#[0m[38;2;145;103;69m9[0m[38;2;156;114;78mB[0m[38;2;156;114;78mB[0m[38;2;155;112;76mB[0m[38;2;159;117;80mB[0m[38;2;167;127;89m&[0m[38;2;177;135;97m&[0m[38;2;179;137;97m&[0m[38;2;178;136;95m&[0m[38;2;178;137;93m&[0m[38;2;178;137;92m&[0m[38;2;178;137;93m&[0m[38;2;179;138;93m&[0m[38;2;178;137;93m&[0m[38;2;176;136;94m&[0m[38;2;166;124;87m&[0m[38;2;143;101;71m9[0m[38;2;116;76;52mG[0m[38;2;97;60;39mM[0m[38;2;101;65;44mH[0m[38;2;112;73;51mG[0m[38;2;117;76;50mG[0m[38;2;128;84;54mS[0m[38;2;130;86;55m#[0m[38;2;133;89;59m#[0m[38;2;137;93;60m#[0m");
	$display("[38;2;81;54;38mh[0m[38;2;101;71;55mG[0m[38;2;129;93;74m#[0m[38;2;150;109;84mB[0m[38;2;160;118;87mB[0m[38;2;162;121;86mB[0m[38;2;162;121;86mB[0m[38;2;162;122;87mB[0m[38;2;162;122;87mB[0m[38;2;162;122;87mB[0m[38;2;164;124;89m&[0m[38;2;165;125;90m&[0m[38;2;166;126;91m&[0m[38;2;161;121;86mB[0m[38;2;152;110;75mB[0m[38;2;146;103;70m9[0m[38;2;144;101;69m9[0m[38;2;144;101;70m9[0m[38;2;147;105;75m9[0m[38;2;132;94;63m#[0m[38;2;125;89;55mS[0m[38;2;152;116;76mB[0m[38;2;178;141;95m&[0m[38;2;181;147;95m&[0m[38;2;151;118;74mB[0m[38;2;132;98;63m#[0m[38;2;125;92;60m#[0m[38;2;111;77;43mG[0m[38;2;145;108;65m9[0m[38;2;149;113;65m9[0m[38;2;151;113;68mB[0m[38;2;150;112;66m9[0m[38;2;150;112;66m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;148;111;65m9[0m[38;2;151;119;79mB[0m[38;2;167;150;111m@[0m[38;2;72;62;44mh[0m[38;2;52;31;21mA[0m[38;2;164;129;100m&[0m[38;2;196;160;113m@[0m[38;2;197;162;109m@[0m[38;2;195;158;115m@[0m[38;2;181;145;107m@[0m[38;2;188;153;114m@[0m[38;2;194;160;116m@[0m[38;2;196;162;115m@[0m[38;2;197;162;115m@[0m[38;2;197;162;116m@[0m[38;2;198;164;117m@[0m[38;2;198;164;115m@[0m[38;2;198;164;118m@[0m[38;2;199;165;120m@[0m[38;2;195;162;116m@[0m[38;2;194;161;116m@[0m[38;2;194;161;117m@[0m[38;2;189;156;112m@[0m[38;2;194;161;116m@[0m[38;2;194;162;116m@[0m[38;2;187;154;112m@[0m[38;2;186;152;111m@[0m[38;2;189;156;113m@[0m[38;2;194;159;118m@[0m[38;2;195;163;121m@[0m[38;2;197;163;114m@[0m[38;2;197;163;115m@[0m[38;2;181;153;115m@[0m[38;2;78;59;37mh[0m[38;2;76;61;43mh[0m[38;2;170;154;118m@[0m[38;2;177;160;121m@[0m[38;2;134;120;93mB[0m[38;2;52;40;23m2[0m[38;2;96;85;74mS[0m[38;2;42;32;18mX[0m[38;2;67;55;43mh[0m[38;2;58;47;35m5[0m[38;2;80;65;49mM[0m[38;2;103;90;71mS[0m[38;2;37;25;17ms[0m[38;2;126;114;86m9[0m[38;2;175;161;125m@[0m[38;2;174;159;121m@[0m[38;2;178;159;121m@[0m[38;2;163;138;104m&[0m[38;2;122;92;55mS[0m[38;2;124;92;52mS[0m[38;2;123;91;50mS[0m[38;2;124;90;50mS[0m[38;2;124;89;48mS[0m[38;2;145;108;66m9[0m[38;2;159;122;78mB[0m[38;2;160;123;78mB[0m[38;2;160;123;79mB[0m[38;2;161;123;79mB[0m[38;2;139;108;69m9[0m[38;2;91;67;35mM[0m[38;2;105;74;46mG[0m[38;2;129;93;60m#[0m[38;2;126;90;55m#[0m[38;2;131;92;57m#[0m[38;2;150;106;70m9[0m[38;2;157;112;77mB[0m[38;2;156;111;76mB[0m[38;2;159;115;79mB[0m[38;2;169;126;88m&[0m[38;2;176;133;95m&[0m[38;2;178;136;96m&[0m[38;2;177;136;95m&[0m[38;2;177;135;95m&[0m[38;2;177;135;95m&[0m[38;2;177;135;94m&[0m[38;2;177;135;94m&[0m[38;2;179;135;97m&[0m[38;2;178;135;95m&[0m[38;2;162;122;85mB[0m[38;2;130;89;64m#[0m[38;2;99;60;43mH[0m[38;2;89;53;36mh[0m[38;2;99;62;39mM[0m[38;2;115;77;49mG[0m[38;2;129;88;58m#[0m[38;2;119;82;51mS[0m[38;2;111;74;44mG[0m[38;2;115;78;50mG[0m[38;2;114;77;50mG[0m[38;2;109;72;47mG[0m[38;2;104;67;45mH[0m");
	$display("[38;2;90;62;42mM[0m[38;2;79;53;38mh[0m[38;2;73;48;37m3[0m[38;2;82;55;41mh[0m[38;2;101;72;53mG[0m[38;2;120;90;65m#[0m[38;2;145;110;79mB[0m[38;2;159;120;86mB[0m[38;2;164;121;87m&[0m[38;2;162;121;86mB[0m[38;2;163;123;88m&[0m[38;2;162;123;88m&[0m[38;2;163;123;88m&[0m[38;2;165;125;90m&[0m[38;2;165;126;91m&[0m[38;2;162;123;87m&[0m[38;2;154;115;79mB[0m[38;2;146;107;72m9[0m[38;2;149;110;72m9[0m[38;2;149;109;74mB[0m[38;2;136;97;68m9[0m[38;2;124;86;58mS[0m[38;2;136;98;68m9[0m[38;2;163;130;88m&[0m[38;2;140;108;68m9[0m[38;2;126;94;59m#[0m[38;2;124;91;58m#[0m[38;2;111;76;43mG[0m[38;2;142;106;66m9[0m[38;2;147;111;66m9[0m[38;2;149;111;68m9[0m[38;2;149;111;66m9[0m[38;2;148;112;65m9[0m[38;2;148;112;66m9[0m[38;2;148;112;66m9[0m[38;2;148;111;65m9[0m[38;2;147;111;65m9[0m[38;2;147;111;65m9[0m[38;2;146;111;65m9[0m[38;2;146;112;65m9[0m[38;2;145;111;64m9[0m[38;2;145;111;62m9[0m[38;2;158;130;87m&[0m[38;2;166;153;116m@[0m[38;2;71;59;46mh[0m[38;2;82;54;40mh[0m[38;2;194;153;114m@[0m[38;2;200;159;118m@[0m[38;2;192;156;113m@[0m[38;2;170;136;98m&[0m[38;2;152;118;90mB[0m[38;2;142;108;81m9[0m[38;2;150;116;85mB[0m[38;2;182;148;110m@[0m[38;2;194;162;114m@[0m[38;2;193;161;114m@[0m[38;2;194;161;116m@[0m[38;2;193;161;114m@[0m[38;2;193;161;115m@[0m[38;2;193;160;116m@[0m[38;2;193;160;117m@[0m[38;2;194;160;114m@[0m[38;2;194;161;112m@[0m[38;2;195;163;115m@[0m[38;2;187;157;115m@[0m[38;2;153;125;91mB[0m[38;2;126;98;70m#[0m[38;2;124;95;69m#[0m[38;2;128;99;70m#[0m[38;2;139;107;78m9[0m[38;2;153;123;91mB[0m[38;2;175;144;104m&[0m[38;2;193;157;113m@[0m[38;2;199;164;123m@[0m[38;2;133;108;78m9[0m[38;2;69;53;32m3[0m[38;2;165;150;115m@[0m[38;2;176;158;122m@[0m[38;2;118;103;81m9[0m[38;2;35;22;9mr[0m[38;2;58;46;36m5[0m[38;2;54;45;33m5[0m[38;2;32;24;15mr[0m[38;2;34;26;17ms[0m[38;2;41;29;20mX[0m[38;2;52;45;34m5[0m[38;2;31;25;20ms[0m[38;2;98;85;62mS[0m[38;2;176;157;124m@[0m[38;2;173;156;120m@[0m[38;2;174;157;122m@[0m[38;2;169;151;118m@[0m[38;2;123;98;62m#[0m[38;2;120;89;51mS[0m[38;2;122;90;50mS[0m[38;2;121;88;47mS[0m[38;2;122;86;45mS[0m[38;2;144;107;66m9[0m[38;2;159;122;78mB[0m[38;2;160;123;78mB[0m[38;2;161;123;79mB[0m[38;2;161;124;80mB[0m[38;2;140;110;70m9[0m[38;2;90;67;37mM[0m[38;2;97;67;43mH[0m[38;2;112;77;49mG[0m[38;2;129;90;60m#[0m[38;2;149;106;72m9[0m[38;2;155;110;72mB[0m[38;2;159;115;78mB[0m[38;2;167;126;89m&[0m[38;2;176;135;95m&[0m[38;2;177;136;96m&[0m[38;2;175;135;94m&[0m[38;2;174;135;93m&[0m[38;2;175;135;94m&[0m[38;2;176;134;95m&[0m[38;2;177;134;93m&[0m[38;2;176;134;93m&[0m[38;2;178;136;96m&[0m[38;2;168;127;92m&[0m[38;2;135;95;68m#[0m[38;2;97;59;40mM[0m[38;2;88;53;36mh[0m[38;2;95;62;43mM[0m[38;2;102;69;46mH[0m[38;2;109;73;48mG[0m[38;2;108;69;45mG[0m[38;2;110;72;50mG[0m[38;2;100;65;42mH[0m[38;2;94;61;39mM[0m[38;2;98;66;44mH[0m[38;2;99;66;42mH[0m[38;2;103;68;41mH[0m[38;2;112;75;44mG[0m");
	$display("[38;2;90;65;43mM[0m[38;2;96;67;45mH[0m[38;2;96;65;45mH[0m[38;2;86;58;43mM[0m[38;2;76;50;38mh[0m[38;2;69;45;34m3[0m[38;2;75;52;39mh[0m[38;2;105;76;59mG[0m[38;2;140;104;81m9[0m[38;2;158;118;87mB[0m[38;2;161;120;86mB[0m[38;2;162;121;86mB[0m[38;2;162;121;86mB[0m[38;2;162;123;87m&[0m[38;2;164;126;90m&[0m[38;2;165;127;91m&[0m[38;2;167;129;93m&[0m[38;2;164;126;90m&[0m[38;2;156;119;83mB[0m[38;2;149;110;74mB[0m[38;2;145;104;71m9[0m[38;2;137;97;68m9[0m[38;2;124;87;61m#[0m[38;2;121;87;58mS[0m[38;2;112;81;51mG[0m[38;2;117;89;58mS[0m[38;2;118;90;57mS[0m[38;2;108;76;42mG[0m[38;2;139;104;64m9[0m[38;2;145;109;63m9[0m[38;2;146;109;65m9[0m[38;2;147;110;64m9[0m[38;2;147;110;64m9[0m[38;2;146;109;65m9[0m[38;2;146;109;64m9[0m[38;2;146;109;64m9[0m[38;2;146;109;64m9[0m[38;2;146;109;64m9[0m[38;2;144;110;64m9[0m[38;2;144;110;64m9[0m[38;2;142;109;63m9[0m[38;2;142;110;62m9[0m[38;2;145;117;80mB[0m[38;2;163;148;116m&[0m[38;2;71;59;43mh[0m[38;2;82;58;41mh[0m[38;2;183;150;113m@[0m[38;2;161;131;96m&[0m[38;2;130;104;76m9[0m[38;2;119;96;70m#[0m[38;2;127;104;78m9[0m[38;2;122;102;73m#[0m[38;2;122;99;73m#[0m[38;2;139;112;82mB[0m[38;2;177;148;108m@[0m[38;2;191;159;114m@[0m[38;2;193;159;114m@[0m[38;2;193;160;115m@[0m[38;2;193;160;115m@[0m[38;2;193;160;115m@[0m[38;2;192;160;116m@[0m[38;2;193;159;115m@[0m[38;2;192;159;115m@[0m[38;2;169;139;99m&[0m[38;2;139;113;78m9[0m[38;2;134;110;78m9[0m[38;2;135;112;81m9[0m[38;2;141;118;87mB[0m[38;2;147;121;89mB[0m[38;2;141;115;83mB[0m[38;2;126;103;73m9[0m[38;2;115;96;68m#[0m[38;2;118;98;71m#[0m[38;2;138;114;86mB[0m[38;2;118;94;71m#[0m[38;2;68;53;36m3[0m[38;2;163;151;115m@[0m[38;2;173;158;119m@[0m[38;2;107;90;66mS[0m[38;2;59;46;34m5[0m[38;2;31;24;16mr[0m[38;2;31;25;12mr[0m[38;2;44;32;20mX[0m[38;2;53;42;27m2[0m[38;2;54;40;25m2[0m[38;2;37;27;17ms[0m[38;2;33;25;14mr[0m[38;2;74;61;43mh[0m[38;2;169;151;121m@[0m[38;2;170;154;116m@[0m[38;2;159;143;108m&[0m[38;2;171;156;121m@[0m[38;2;132;112;74m9[0m[38;2;117;87;49mS[0m[38;2;120;88;47mS[0m[38;2;119;88;44mS[0m[38;2;121;85;44mS[0m[38;2;143;105;64m9[0m[38;2;160;122;79mB[0m[38;2;161;123;79mB[0m[38;2;162;123;80mB[0m[38;2;162;124;81mB[0m[38;2;140;110;71m9[0m[38;2;87;62;36mM[0m[38;2;98;65;44mH[0m[38;2;125;89;61m#[0m[38;2;143;103;70m9[0m[38;2;157;113;78mB[0m[38;2;171;126;89m&[0m[38;2;176;134;96m&[0m[38;2;175;136;98m&[0m[38;2;174;136;96m&[0m[38;2;174;135;94m&[0m[38;2;174;135;94m&[0m[38;2;174;135;93m&[0m[38;2;175;134;94m&[0m[38;2;176;134;93m&[0m[38;2;176;134;92m&[0m[38;2;176;134;96m&[0m[38;2;151;111;80mB[0m[38;2;122;83;61mS[0m[38;2;102;64;45mH[0m[38;2;94;60;41mM[0m[38;2;99;68;47mH[0m[38;2;91;63;39mM[0m[38;2;82;54;31mh[0m[38;2;85;54;35mh[0m[38;2;91;58;40mM[0m[38;2;100;66;46mH[0m[38;2;99;65;42mH[0m[38;2;99;64;38mH[0m[38;2;117;81;49mS[0m[38;2;133;97;57m#[0m[38;2;149;112;67m9[0m[38;2;161;123;75mB[0m");
	$display("[38;2;65;45;27m5[0m[38;2;69;45;29m5[0m[38;2;79;51;34mh[0m[38;2;87;59;40mM[0m[38;2;92;65;44mH[0m[38;2;91;64;46mH[0m[38;2;82;58;42mM[0m[38;2;72;48;34m3[0m[38;2;74;49;34m3[0m[38;2;105;75;57mG[0m[38;2;143;108;84mB[0m[38;2;159;118;86mB[0m[38;2;159;118;82mB[0m[38;2;159;121;84mB[0m[38;2;160;123;87mB[0m[38;2;162;124;88m&[0m[38;2;163;126;90m&[0m[38;2;166;128;92m&[0m[38;2;166;128;93m&[0m[38;2;164;125;90m&[0m[38;2;157;117;82mB[0m[38;2;148;109;77mB[0m[38;2;138;102;72m9[0m[38;2;127;92;64m#[0m[38;2;103;71;46mH[0m[38;2;101;73;49mG[0m[38;2;105;79;51mG[0m[38;2;105;75;42mG[0m[38;2;139;104;60m9[0m[38;2;144;109;61m9[0m[38;2;145;108;64m9[0m[38;2;145;108;64m9[0m[38;2;145;108;64m9[0m[38;2;145;108;64m9[0m[38;2;144;108;63m9[0m[38;2;144;107;63m9[0m[38;2;144;107;63m9[0m[38;2;144;107;63m9[0m[38;2;142;108;63m9[0m[38;2;142;108;63m9[0m[38;2;140;107;61m9[0m[38;2;138;108;62m9[0m[38;2;139;113;77m9[0m[38;2;162;147;112m&[0m[38;2;72;63;45mh[0m[38;2;77;59;46mM[0m[38;2;122;98;71m#[0m[38;2;120;96;65m#[0m[38;2;153;127;92m&[0m[38;2;176;147;108m@[0m[38;2;186;153;111m@[0m[38;2;189;153;113m@[0m[38;2;184;150;111m@[0m[38;2;169;139;98m&[0m[38;2;174;146;103m&[0m[38;2;188;157;112m@[0m[38;2;192;158;113m@[0m[38;2;192;159;114m@[0m[38;2;191;158;113m@[0m[38;2;191;158;113m@[0m[38;2;191;159;115m@[0m[38;2;191;158;115m@[0m[38;2;189;156;116m@[0m[38;2;174;142;103m&[0m[38;2;178;145;107m@[0m[38;2;189;154;114m@[0m[38;2;192;159;115m@[0m[38;2;195;160;116m@[0m[38;2;196;156;115m@[0m[38;2;196;156;114m@[0m[38;2;192;154;112m@[0m[38;2;182;148;108m@[0m[38;2;164;134;98m&[0m[38;2;137;109;78m9[0m[38;2;88;68;47mH[0m[38;2;69;57;42mh[0m[38;2;165;151;119m@[0m[38;2;166;148;113m&[0m[38;2;101;80;58mG[0m[38;2;103;82;66mS[0m[38;2;64;43;24m5[0m[38;2;122;97;72m#[0m[38;2;138;104;84m9[0m[38;2;124;91;74m#[0m[38;2;112;87;63mS[0m[38;2;116;90;72m#[0m[38;2;49;30;19mX[0m[38;2;51;43;25m2[0m[38;2;155;140;111m&[0m[38;2;169;155;117m@[0m[38;2;155;140;103m&[0m[38;2;171;155;118m@[0m[38;2;146;127;90mB[0m[38;2;114;85;49mS[0m[38;2;118;86;47mS[0m[38;2;116;86;45mS[0m[38;2;119;84;44mS[0m[38;2;143;105;61m9[0m[38;2;158;121;76mB[0m[38;2;159;123;78mB[0m[38;2;158;123;80mB[0m[38;2;147;111;71m9[0m[38;2;120;88;53mS[0m[38;2;100;68;44mH[0m[38;2;124;83;60mS[0m[38;2;150;107;76mB[0m[38;2;167;123;88m&[0m[38;2;177;132;95m&[0m[38;2;176;134;95m&[0m[38;2;174;134;95m&[0m[38;2;174;134;98m&[0m[38;2;174;134;97m&[0m[38;2;173;134;95m&[0m[38;2;173;135;95m&[0m[38;2;174;135;94m&[0m[38;2;175;133;93m&[0m[38;2;174;134;95m&[0m[38;2;165;130;93m&[0m[38;2;126;92;65m#[0m[38;2;92;57;40mM[0m[38;2;95;61;46mH[0m[38;2;96;65;44mH[0m[38;2;92;63;38mM[0m[38;2;81;54;31mh[0m[38;2;77;50;29m3[0m[38;2;80;53;32mh[0m[38;2;92;61;38mM[0m[38;2;106;73;45mG[0m[38;2;133;98;63m#[0m[38;2;138;102;65m9[0m[38;2;141;104;62m9[0m[38;2;161;124;76mB[0m[38;2;167;128;76mB[0m[38;2;166;126;74mB[0m[38;2;164;126;74mB[0m");
	$display("[38;2;72;52;34m3[0m[38;2;67;48;32m3[0m[38;2;62;42;27m5[0m[38;2;60;38;24m2[0m[38;2;63;40;25m2[0m[38;2;71;47;31m3[0m[38;2;83;56;40mh[0m[38;2;91;64;50mH[0m[38;2;82;58;46mM[0m[38;2;71;48;35m3[0m[38;2;84;57;41mM[0m[38;2;118;85;64mS[0m[38;2;152;115;84mB[0m[38;2;159;119;83mB[0m[38;2;159;119;83mB[0m[38;2;159;120;84mB[0m[38;2;160;123;87mB[0m[38;2;163;124;88m&[0m[38;2;164;126;91m&[0m[38;2;165;127;91m&[0m[38;2;165;127;90m&[0m[38;2;163;125;89m&[0m[38;2;158;120;87mB[0m[38;2;150;112;82mB[0m[38;2;126;90;65m#[0m[38;2;107;74;53mG[0m[38;2;96;66;43mH[0m[38;2;99;69;40mH[0m[38;2;133;98;61m#[0m[38;2;143;107;63m9[0m[38;2;144;106;64m9[0m[38;2;142;106;64m9[0m[38;2;142;106;61m9[0m[38;2;142;106;61m9[0m[38;2;141;105;63m9[0m[38;2;140;105;62m9[0m[38;2;139;105;60m9[0m[38;2;140;105;60m9[0m[38;2;139;105;60m9[0m[38;2;139;105;60m9[0m[38;2;139;106;60m9[0m[38;2;137;105;61m9[0m[38;2;122;104;68m#[0m[38;2;159;146;112m&[0m[38;2;75;64;46mM[0m[38;2;60;43;28m5[0m[38;2;158;127;93m&[0m[38;2;188;148;108m@[0m[38;2;193;151;110m@[0m[38;2;191;149;110m@[0m[38;2;192;150;109m@[0m[38;2;192;154;113m@[0m[38;2;193;156;114m@[0m[38;2;194;158;116m@[0m[38;2;191;156;114m@[0m[38;2;192;158;116m@[0m[38;2;161;128;89m&[0m[38;2;156;122;86mB[0m[38;2;190;157;118m@[0m[38;2;190;157;114m@[0m[38;2;190;157;113m@[0m[38;2;190;157;114m@[0m[38;2;190;157;114m@[0m[38;2;192;158;115m@[0m[38;2;192;158;115m@[0m[38;2;190;156;114m@[0m[38;2;189;153;111m@[0m[38;2;189;149;108m@[0m[38;2;189;146;107m@[0m[38;2;191;145;108m@[0m[38;2;191;145;106m@[0m[38;2;193;149;108m@[0m[38;2;192;151;109m@[0m[38;2;194;153;114m@[0m[38;2;122;94;71m#[0m[38;2;78;64;45mM[0m[38;2;171;151;121m@[0m[38;2;147;130;104m&[0m[38;2;91;71;49mH[0m[38;2;112;85;63mS[0m[38;2;140;109;87mB[0m[38;2;100;73;59mG[0m[38;2;62;35;26m2[0m[38;2;45;24;19mX[0m[38;2;43;22;17ms[0m[38;2;112;78;66mS[0m[38;2;88;64;50mH[0m[38;2;33;28;13ms[0m[38;2;137;123;96mB[0m[38;2;173;156;119m@[0m[38;2;155;140;103m&[0m[38;2;169;152;117m@[0m[38;2;158;140;104m&[0m[38;2;112;88;51mS[0m[38;2;115;84;45mG[0m[38;2;116;83;43mG[0m[38;2;115;83;42mG[0m[38;2;133;101;61m#[0m[38;2;155;121;79mB[0m[38;2;147;113;69m9[0m[38;2;130;97;60m#[0m[38;2;120;86;59mS[0m[38;2;125;90;62m#[0m[38;2;137;101;67m9[0m[38;2;163;123;85mB[0m[38;2;174;132;95m&[0m[38;2;176;132;93m&[0m[38;2;175;133;93m&[0m[38;2;173;134;95m&[0m[38;2;172;133;95m&[0m[38;2;173;133;96m&[0m[38;2;173;132;94m&[0m[38;2;171;134;92m&[0m[38;2;171;134;93m&[0m[38;2;173;132;95m&[0m[38;2;173;132;97m&[0m[38;2;151;114;82mB[0m[38;2;110;76;50mG[0m[38;2;98;66;43mH[0m[38;2;106;74;51mG[0m[38;2;95;64;42mH[0m[38;2;86;56;34mh[0m[38;2;81;52;30m3[0m[38;2;82;55;32mh[0m[38;2;87;59;36mM[0m[38;2;99;67;42mH[0m[38;2;125;89;58m#[0m[38;2;145;106;68m9[0m[38;2;165;125;81mB[0m[38;2;160;123;77mB[0m[38;2;161;124;78mB[0m[38;2;170;132;84m&[0m[38;2;169;131;82m&[0m[38;2;167;128;78m&[0m[38;2;162;125;75mB[0m");
	$display("[38;2;117;90;52mS[0m[38;2;106;80;46mG[0m[38;2;94;69;41mH[0m[38;2;82;58;35mh[0m[38;2;72;50;30m3[0m[38;2;67;43;27m5[0m[38;2;62;39;24m2[0m[38;2;67;43;28m5[0m[38;2;79;53;38mh[0m[38;2;87;60;43mM[0m[38;2;80;56;40mh[0m[38;2;72;48;34m3[0m[38;2;96;65;48mH[0m[38;2;139;100;77m9[0m[38;2;157;117;85mB[0m[38;2;159;118;83mB[0m[38;2;159;119;83mB[0m[38;2;159;121;86mB[0m[38;2;160;121;87mB[0m[38;2;163;125;87m&[0m[38;2;165;126;87m&[0m[38;2;164;125;88m&[0m[38;2;164;125;90m&[0m[38;2;164;125;91m&[0m[38;2;159;119;89mB[0m[38;2;148;108;83mB[0m[38;2;122;87;62m#[0m[38;2;101;69;44mH[0m[38;2;107;75;46mG[0m[38;2;121;87;51mS[0m[38;2;135;99;62m#[0m[38;2;138;106;62m9[0m[38;2;136;105;59m9[0m[38;2;137;104;59m9[0m[38;2;139;103;59m9[0m[38;2;138;103;58m9[0m[38;2;136;104;58m#[0m[38;2;136;103;58m#[0m[38;2;136;103;58m#[0m[38;2;136;103;60m9[0m[38;2;136;103;60m9[0m[38;2;129;98;59m#[0m[38;2;97;82;51mG[0m[38;2;158;144;112m&[0m[38;2;81;69;53mH[0m[38;2;42;27;11ms[0m[38;2;161;123;93m&[0m[38;2;192;142;104m@[0m[38;2;192;140;101m@[0m[38;2;189;139;103m@[0m[38;2;192;142;104m@[0m[38;2;193;148;109m@[0m[38;2;193;154;112m@[0m[38;2;191;157;114m@[0m[38;2;189;156;113m@[0m[38;2;189;156;115m@[0m[38;2;175;142;103m&[0m[38;2;183;149;111m@[0m[38;2;189;156;116m@[0m[38;2;189;156;114m@[0m[38;2;189;156;113m@[0m[38;2;189;156;113m@[0m[38;2;189;156;113m@[0m[38;2;190;157;114m@[0m[38;2;190;156;113m@[0m[38;2;190;153;111m@[0m[38;2;189;147;107m@[0m[38;2;189;142;104m@[0m[38;2;190;140;102m@[0m[38;2;191;139;104m@[0m[38;2;190;139;102m@[0m[38;2;191;141;102m@[0m[38;2;190;140;103m@[0m[38;2;193;143;108m@[0m[38;2;114;83;62mS[0m[38;2;88;75;54mH[0m[38;2;172;154;123m@[0m[38;2;118;101;80m9[0m[38;2;103;78;49mG[0m[38;2;173;142;110m&[0m[38;2;95;67;50mH[0m[38;2;40;21;18ms[0m[38;2;43;27;24mX[0m[38;2;42;22;17ms[0m[38;2;53;25;19mX[0m[38;2;132;100;80m9[0m[38;2;84;64;45mM[0m[38;2;30;20;13mr[0m[38;2;116;100;80m#[0m[38;2;173;155;121m@[0m[38;2;155;140;106m&[0m[38;2;163;146;115m&[0m[38;2;168;150;118m@[0m[38;2;118;98;60m#[0m[38;2;111;85;43mG[0m[38;2;111;83;47mG[0m[38;2;103;77;49mG[0m[38;2;81;60;37mh[0m[38;2;91;68;49mH[0m[38;2;111;83;57mS[0m[38;2;126;90;57m#[0m[38;2;147;107;74m9[0m[38;2;164;125;88m&[0m[38;2;173;134;95m&[0m[38;2;173;134;94m&[0m[38;2;172;133;94m&[0m[38;2;172;133;94m&[0m[38;2;172;133;94m&[0m[38;2;172;133;94m&[0m[38;2;172;132;93m&[0m[38;2;172;131;91m&[0m[38;2;172;132;91m&[0m[38;2;173;132;91m&[0m[38;2;173;134;96m&[0m[38;2;164;125;92m&[0m[38;2;130;94;65m#[0m[38;2;105;69;44mH[0m[38;2;112;76;52mG[0m[38;2;116;80;56mS[0m[38;2;102;68;42mH[0m[38;2;83;55;30mh[0m[38;2;85;56;33mh[0m[38;2;95;66;42mH[0m[38;2;103;74;47mG[0m[38;2;107;78;48mG[0m[38;2;111;80;46mG[0m[38;2;132;95;59m#[0m[38;2;145;103;64m9[0m[38;2;151;109;66m9[0m[38;2;149;109;66m9[0m[38;2;147;108;65m9[0m[38;2;150;111;68m9[0m[38;2;160;121;77mB[0m[38;2;167;130;83m&[0m[38;2;168;130;82m&[0m");
	$display("[38;2;136;103;58m#[0m[38;2;136;103;59m#[0m[38;2;134;102;60m#[0m[38;2;130;98;58m#[0m[38;2;123;91;54mS[0m[38;2;110;81;47mG[0m[38;2;96;69;39mH[0m[38;2;80;56;32mh[0m[38;2;69;47;29m5[0m[38;2;65;44;28m5[0m[38;2;73;52;33m3[0m[38;2;84;61;39mM[0m[38;2;84;58;37mh[0m[38;2;84;56;38mh[0m[38;2;109;79;58mS[0m[38;2;143;109;82mB[0m[38;2;156;117;86mB[0m[38;2;159;116;82mB[0m[38;2;159;117;83mB[0m[38;2;159;120;86mB[0m[38;2;162;122;88m&[0m[38;2;164;124;91m&[0m[38;2;165;125;93m&[0m[38;2;165;125;91m&[0m[38;2;165;123;90m&[0m[38;2;167;124;92m&[0m[38;2;161;122;89m&[0m[38;2;145;109;77m9[0m[38;2;126;90;59m#[0m[38;2;112;77;49mG[0m[38;2;93;67;48mH[0m[38;2;82;61;40mM[0m[38;2;84;64;37mM[0m[38;2;107;83;51mG[0m[38;2;128;98;59m#[0m[38;2;137;103;60m9[0m[38;2;138;102;58m#[0m[38;2;134;101;57m#[0m[38;2;133;101;56m#[0m[38;2;133;101;58m#[0m[38;2;134;101;60m#[0m[38;2;127;94;60m#[0m[38;2;84;67;46mM[0m[38;2;153;136;111m&[0m[38;2;90;80;62mG[0m[38;2;26;19;8mi[0m[38;2;121;88;67m#[0m[38;2;189;142;107m@[0m[38;2;192;141;103m@[0m[38;2;189;143;107m@[0m[38;2;191;147;108m@[0m[38;2;191;152;111m@[0m[38;2;190;156;113m@[0m[38;2;189;157;113m@[0m[38;2;189;156;113m@[0m[38;2;189;156;113m@[0m[38;2;190;157;114m@[0m[38;2;190;157;112m@[0m[38;2;189;157;112m@[0m[38;2;189;157;112m@[0m[38;2;189;157;112m@[0m[38;2;189;156;113m@[0m[38;2;189;156;114m@[0m[38;2;189;156;115m@[0m[38;2;190;156;114m@[0m[38;2;190;154;113m@[0m[38;2;190;152;111m@[0m[38;2;191;150;109m@[0m[38;2;191;147;108m@[0m[38;2;190;146;107m@[0m[38;2;190;146;106m@[0m[38;2;190;145;105m@[0m[38;2;191;146;106m@[0m[38;2;192;148;112m@[0m[38;2;99;74;52mG[0m[38;2;100;89;66mS[0m[38;2;169;152;121m@[0m[38;2;86;67;51mH[0m[38;2;114;83;69mS[0m[38;2;129;98;82m9[0m[38;2;64;40;30m5[0m[38;2;40;21;16ms[0m[38;2;52;29;23mA[0m[38;2;89;60;43mM[0m[38;2;142;110;83mB[0m[38;2;124;98;75m#[0m[38;2;43;28;17mX[0m[38;2;30;20;14mr[0m[38;2;86;73;55mH[0m[38;2;169;152;120m@[0m[38;2;156;139;105m&[0m[38;2;150;132;104m&[0m[38;2;173;155;122m@[0m[38;2;135;114;82m9[0m[38;2;91;68;42mH[0m[38;2;85;64;41mM[0m[38;2;88;71;48mH[0m[38;2;60;48;33m5[0m[38;2;27;16;9mi[0m[38;2;68;46;33m3[0m[38;2;157;119;88mB[0m[38;2;174;131;91m&[0m[38;2;173;132;93m&[0m[38;2;172;131;94m&[0m[38;2;171;131;95m&[0m[38;2;170;132;96m&[0m[38;2;171;132;95m&[0m[38;2;171;132;94m&[0m[38;2;171;132;93m&[0m[38;2;172;131;92m&[0m[38;2;172;132;92m&[0m[38;2;173;132;94m&[0m[38;2;171;130;95m&[0m[38;2;146;106;77m9[0m[38;2;111;75;49mG[0m[38;2;105;72;49mG[0m[38;2;112;79;56mS[0m[38;2;107;74;51mG[0m[38;2;101;69;43mH[0m[38;2;107;76;48mG[0m[38;2;101;71;43mH[0m[38;2;105;75;49mG[0m[38;2;107;77;50mG[0m[38;2;107;77;47mG[0m[38;2;106;76;45mG[0m[38;2;107;76;45mG[0m[38;2;125;91;56m#[0m[38;2;137;100;60m#[0m[38;2;152;112;68mB[0m[38;2;159;118;73mB[0m[38;2;157;119;73mB[0m[38;2;149;113;68m9[0m[38;2;143;106;61m9[0m[38;2;147;110;65m9[0m[38;2;159;121;75mB[0m");
	$display("[38;2;133;100;59m#[0m[38;2;134;101;58m#[0m[38;2;134;101;58m#[0m[38;2;133;100;60m#[0m[38;2;134;100;61m#[0m[38;2;135;102;60m#[0m[38;2;134;101;59m#[0m[38;2;129;97;59m#[0m[38;2;116;87;53mS[0m[38;2;99;72;41mH[0m[38;2;79;54;30m3[0m[38;2;68;45;29m5[0m[38;2;73;49;36m3[0m[38;2;81;56;41mh[0m[38;2;82;54;38mh[0m[38;2;88;60;43mM[0m[38;2;118;86;65mS[0m[38;2;150;112;84mB[0m[38;2;160;118;86mB[0m[38;2;159;116;83mB[0m[38;2;159;118;84mB[0m[38;2;161;120;87mB[0m[38;2;162;122;90m&[0m[38;2;163;123;91m&[0m[38;2;165;125;92m&[0m[38;2;165;125;93m&[0m[38;2;164;125;92m&[0m[38;2;166;127;93m&[0m[38;2;157;122;93m&[0m[38;2;84;65;49mM[0m[38;2;21;15;9m;[0m[38;2;31;22;12mr[0m[38;2;65;50;38m3[0m[38;2;80;66;51mM[0m[38;2;84;68;45mM[0m[38;2;92;70;40mH[0m[38;2;118;90;57mS[0m[38;2;131;100;60m#[0m[38;2;132;100;56m#[0m[38;2;132;99;55m#[0m[38;2;133;99;58m#[0m[38;2;128;97;60m#[0m[38;2;81;67;45mM[0m[38;2;145;130;106m&[0m[38;2;100;91;68mS[0m[38;2;22;19;11mi[0m[38;2;72;51;34m3[0m[38;2;180;145;106m@[0m[38;2;191;152;109m@[0m[38;2;190;154;114m@[0m[38;2;189;155;110m@[0m[38;2;189;154;112m@[0m[38;2;189;155;112m@[0m[38;2;188;156;113m@[0m[38;2;189;156;113m@[0m[38;2;189;156;112m@[0m[38;2;192;159;115m@[0m[38;2;190;158;114m@[0m[38;2;190;157;112m@[0m[38;2;191;157;111m@[0m[38;2;192;157;114m@[0m[38;2;192;159;112m@[0m[38;2;193;160;114m@[0m[38;2;189;157;115m@[0m[38;2;188;155;116m@[0m[38;2;187;155;114m@[0m[38;2;186;156;113m@[0m[38;2;187;156;112m@[0m[38;2;190;155;113m@[0m[38;2;189;155;110m@[0m[38;2;190;154;111m@[0m[38;2;191;154;112m@[0m[38;2;190;154;112m@[0m[38;2;186;152;114m@[0m[38;2;83;65;42mM[0m[38;2;118;109;82m9[0m[38;2;153;136;107m&[0m[38;2;63;45;31m5[0m[38;2;108;81;67mS[0m[38;2;93;66;51mH[0m[38;2;97;69;49mH[0m[38;2;120;90;66m#[0m[38;2;135;104;79m9[0m[38;2;130;102;76m9[0m[38;2;84;63;51mM[0m[38;2;36;24;18ms[0m[38;2;32;22;13mr[0m[38;2;32;21;14mr[0m[38;2;57;46;32m5[0m[38;2;157;143;109m&[0m[38;2;161;145;107m&[0m[38;2;123;107;82m9[0m[38;2;140;124;103mB[0m[38;2;89;75;56mH[0m[38;2;52;42;29m2[0m[38;2;39;32;20mX[0m[38;2;48;39;25mA[0m[38;2;64;48;33m5[0m[38;2;54;45;28m2[0m[38;2;32;19;7mi[0m[38;2;117;86;68m#[0m[38;2;172;131;98m&[0m[38;2;171;131;94m&[0m[38;2;171;131;95m&[0m[38;2;171;131;95m&[0m[38;2;171;131;95m&[0m[38;2;171;131;96m&[0m[38;2;171;131;94m&[0m[38;2;171;132;92m&[0m[38;2;172;132;94m&[0m[38;2;172;131;97m&[0m[38;2;153;115;87mB[0m[38;2;120;84;61mS[0m[38;2;103;69;50mG[0m[38;2;105;72;52mG[0m[38;2;101;71;48mH[0m[38;2;99;68;43mH[0m[38;2;115;81;53mS[0m[38;2;140;105;71m9[0m[38;2;145;109;72m9[0m[38;2;112;79;47mG[0m[38;2;107;76;47mG[0m[38;2;104;75;47mG[0m[38;2;104;76;45mG[0m[38;2;104;74;43mH[0m[38;2;103;73;43mH[0m[38;2;118;86;53mS[0m[38;2;130;95;56m#[0m[38;2;147;109;63m9[0m[38;2;157;116;69mB[0m[38;2;156;118;71mB[0m[38;2;155;119;72mB[0m[38;2;154;118;72mB[0m[38;2;144;106;62m9[0m[38;2;139;100;57m#[0m");
	$display("[38;2;132;98;59m#[0m[38;2;132;99;58m#[0m[38;2;132;99;58m#[0m[38;2;132;98;60m#[0m[38;2;132;98;60m#[0m[38;2;133;99;58m#[0m[38;2;132;100;58m#[0m[38;2;133;100;58m#[0m[38;2;134;100;59m#[0m[38;2;136;99;60m#[0m[38;2;128;95;57m#[0m[38;2;108;83;48mG[0m[38;2;86;64;38mM[0m[38;2;68;45;27m5[0m[38;2;64;40;24m2[0m[38;2;66;45;33m5[0m[38;2;72;49;37m3[0m[38;2;92;61;45mM[0m[38;2;130;92;69m#[0m[38;2;153;113;84mB[0m[38;2;158;118;84mB[0m[38;2;157;117;83mB[0m[38;2;160;118;89mB[0m[38;2;159;120;88mB[0m[38;2;162;125;91m&[0m[38;2;162;127;92m&[0m[38;2;162;128;93m&[0m[38;2;160;127;95m&[0m[38;2;96;73;55mG[0m[38;2;27;19;10mi[0m[38;2;45;36;23mA[0m[38;2;50;38;28m2[0m[38;2;44;35;28mA[0m[38;2;25;21;15mr[0m[38;2;29;28;22ms[0m[38;2;44;39;26mA[0m[38;2;59;46;27m5[0m[38;2;84;65;40mM[0m[38;2;113;88;54mS[0m[38;2;130;98;57m#[0m[38;2;132;98;56m#[0m[38;2;130;99;60m#[0m[38;2;87;69;46mH[0m[38;2;126;109;85m9[0m[38;2;112;100;79m#[0m[38;2;26;19;14mi[0m[38;2;34;21;12mr[0m[38;2;130;105;74m9[0m[38;2;190;157;115m@[0m[38;2;186;155;113m@[0m[38;2;187;155;111m@[0m[38;2;189;154;111m@[0m[38;2;188;154;112m@[0m[38;2;188;155;112m@[0m[38;2;188;155;111m@[0m[38;2;173;138;105m&[0m[38;2;121;89;68m#[0m[38;2;130;104;85m9[0m[38;2;133;106;89m9[0m[38;2;132;103;84m9[0m[38;2;127;99;82m9[0m[38;2;104;79;64mS[0m[38;2;107;80;60mS[0m[38;2;171;139;104m&[0m[38;2;189;155;113m@[0m[38;2;188;155;114m@[0m[38;2;186;156;113m@[0m[38;2;187;156;112m@[0m[38;2;188;155;112m@[0m[38;2;188;155;110m@[0m[38;2;189;154;112m@[0m[38;2;190;154;112m@[0m[38;2;189;155;112m@[0m[38;2;178;146;109m@[0m[38;2;73;55;34m3[0m[38;2;139;129;100mB[0m[38;2;130;109;89m9[0m[38;2;60;36;27m2[0m[38;2;129;90;70m#[0m[38;2;147;108;85mB[0m[38;2;126;100;77m9[0m[38;2;77;63;46mM[0m[38;2;43;35;25mA[0m[38;2;26;22;16mr[0m[38;2;25;20;17mr[0m[38;2;28;24;14mr[0m[38;2;30;24;14mr[0m[38;2;31;21;18mr[0m[38;2;37;26;16ms[0m[38;2;130;116;95mB[0m[38;2;146;132;108m&[0m[38;2;78;66;49mM[0m[38;2;54;42;30m2[0m[38;2;37;28;19ms[0m[38;2;24;19;14mi[0m[38;2;17;13;8m;[0m[38;2;18;13;6m;[0m[38;2;54;42;31m2[0m[38;2;82;65;44mM[0m[38;2;43;30;20mX[0m[38;2;50;32;25mA[0m[38;2;155;121;95mB[0m[38;2;170;130;94m&[0m[38;2;170;130;94m&[0m[38;2;170;130;93m&[0m[38;2;170;131;92m&[0m[38;2;171;131;92m&[0m[38;2;171;132;90m&[0m[38;2;170;133;92m&[0m[38;2;161;124;92m&[0m[38;2;128;91;66m#[0m[38;2;103;68;47mH[0m[38;2;96;66;48mH[0m[38;2;90;64;44mM[0m[38;2;92;65;39mM[0m[38;2;112;83;48mG[0m[38;2;138;105;66m9[0m[38;2;154;117;76mB[0m[38;2;154;117;74mB[0m[38;2;143;110;67m9[0m[38;2;109;79;44mG[0m[38;2;103;76;44mG[0m[38;2;102;75;46mG[0m[38;2;103;73;45mH[0m[38;2;102;72;42mH[0m[38;2;103;70;39mH[0m[38;2;116;79;47mG[0m[38;2;125;84;50mS[0m[38;2;138;99;58m#[0m[38;2;149;107;64m9[0m[38;2;149;108;65m9[0m[38;2;148;109;65m9[0m[38;2;146;107;65m9[0m[38;2;145;105;63m9[0m[38;2;140;101;61m9[0m");
	$display("[38;2;131;97;59m#[0m[38;2;131;97;59m#[0m[38;2;131;97;59m#[0m[38;2;131;97;59m#[0m[38;2;132;98;60m#[0m[38;2;132;97;59m#[0m[38;2;132;97;59m#[0m[38;2;132;98;60m#[0m[38;2;132;98;60m#[0m[38;2;134;97;61m#[0m[38;2;132;97;58m#[0m[38;2;131;99;56m#[0m[38;2;128;98;59m#[0m[38;2;117;86;54mS[0m[38;2;93;66;39mM[0m[38;2;65;45;25m5[0m[38;2;53;36;21mA[0m[38;2;57;35;23m2[0m[38;2;70;43;29m5[0m[38;2;96;67;47mH[0m[38;2;133;99;73m9[0m[38;2;156;118;86mB[0m[38;2;160;118;85mB[0m[38;2;157;118;83mB[0m[38;2;157;121;86mB[0m[38;2;161;122;86mB[0m[38;2;160;125;91m&[0m[38;2;122;98;73m#[0m[38;2;48;38;22mA[0m[38;2;71;60;42mh[0m[38;2;88;73;45mH[0m[38;2;52;42;26m2[0m[38;2;19;15;10m;[0m[38;2;12;10;7m:[0m[38;2;10;10;8m:[0m[38;2;16;15;10m;[0m[38;2;30;26;18ms[0m[38;2;46;35;26mA[0m[38;2;59;45;31m5[0m[38;2;77;58;36mh[0m[38;2;105;79;49mG[0m[38;2;126;97;61m#[0m[38;2;105;83;55mG[0m[38;2;95;82;60mG[0m[38;2;117;106;85m9[0m[38;2;30;21;13mr[0m[38;2;26;20;14mr[0m[38;2;49;32;21mA[0m[38;2;150;121;91mB[0m[38;2;190;158;112m@[0m[38;2;188;156;109m@[0m[38;2;188;155;109m@[0m[38;2;188;155;110m@[0m[38;2;188;155;111m@[0m[38;2;188;155;113m@[0m[38;2;163;130;99m&[0m[38;2;45;20;13ms[0m[38;2;31;9;7mi[0m[38;2;54;25;20mX[0m[38;2;64;28;29m2[0m[38;2;64;28;27m2[0m[38;2;46;18;17ms[0m[38;2;58;31;22mA[0m[38;2;164;131;100m&[0m[38;2;191;154;112m@[0m[38;2;188;155;113m@[0m[38;2;188;155;113m@[0m[38;2;188;155;111m@[0m[38;2;188;155;111m@[0m[38;2;188;156;109m@[0m[38;2;189;154;114m@[0m[38;2;189;156;110m@[0m[38;2;190;160;112m@[0m[38;2;156;129;99m&[0m[38;2;74;59;38mh[0m[38;2;156;139;114m&[0m[38;2;90;76;59mG[0m[38;2;36;20;12mr[0m[38;2;51;27;21mX[0m[38;2;39;20;14ms[0m[38;2;24;21;12mi[0m[38;2;19;22;14mi[0m[38;2;23;23;18mr[0m[38;2;26;23;19mr[0m[38;2;27;23;18mr[0m[38;2;27;23;15mr[0m[38;2;36;33;23mX[0m[38;2;34;31;19ms[0m[38;2;31;21;11mr[0m[38;2;67;54;44mh[0m[38;2;62;50;41m3[0m[38;2;37;30;21mX[0m[38;2;22;17;10mi[0m[38;2;16;12;5m:[0m[38;2;16;13;6m;[0m[38;2;16;13;6m;[0m[38;2;14;13;5m:[0m[38;2;26;23;17mr[0m[38;2;37;27;19ms[0m[38;2;41;32;22mX[0m[38;2;23;10;9m;[0m[38;2;112;88;66mS[0m[38;2;168;131;93m&[0m[38;2;170;129;89m&[0m[38;2;168;130;93m&[0m[38;2;170;128;92m&[0m[38;2;171;130;95m&[0m[38;2;167;128;95m&[0m[38;2;143;107;78m9[0m[38;2;108;74;51mG[0m[38;2;96;65;44mH[0m[38;2;87;61;39mM[0m[38;2;83;60;37mh[0m[38;2;104;78;51mG[0m[38;2;133;102;67m9[0m[38;2;150;115;73mB[0m[38;2;153;115;72mB[0m[38;2;153;115;73mB[0m[38;2;152;115;73mB[0m[38;2;143;109;67m9[0m[38;2;106;78;44mG[0m[38;2;99;73;43mH[0m[38;2;100;72;45mH[0m[38;2;103;72;42mH[0m[38;2;111;78;44mG[0m[38;2;127;91;54m#[0m[38;2;136;97;61m#[0m[38;2;138;97;60m#[0m[38;2;137;98;58m#[0m[38;2;140;99;58m#[0m[38;2;140;99;57m#[0m[38;2;139;99;57m#[0m[38;2;138;98;56m#[0m[38;2;138;97;56m#[0m[38;2;139;98;59m#[0m");
	$display("[38;2;129;95;57m#[0m[38;2;129;95;57m#[0m[38;2;129;95;57m#[0m[38;2;129;96;57m#[0m[38;2;130;96;58m#[0m[38;2;130;96;58m#[0m[38;2;130;96;58m#[0m[38;2;130;96;58m#[0m[38;2;129;96;58m#[0m[38;2;130;96;58m#[0m[38;2;130;96;57m#[0m[38;2;130;96;55m#[0m[38;2;131;96;55m#[0m[38;2;131;97;56m#[0m[38;2;129;96;58m#[0m[38;2;118;90;55mS[0m[38;2;92;70;43mH[0m[38;2;62;43;25m5[0m[38;2;49;31;18mX[0m[38;2;54;34;23mA[0m[38;2;71;47;36m3[0m[38;2;104;71;55mG[0m[38;2;140;100;77m9[0m[38;2;157;117;84mB[0m[38;2;159;119;83mB[0m[38;2;161;117;82mB[0m[38;2;150;115;91mB[0m[38;2;54;39;28m2[0m[38;2;26;22;13mr[0m[38;2;48;37;26mA[0m[38;2;47;40;26mA[0m[38;2;31;26;19ms[0m[38;2;32;25;18ms[0m[38;2;29;24;17mr[0m[38;2;20;18;14mi[0m[38;2;13;12;9m:[0m[38;2;12;10;7m:[0m[38;2;17;12;9m;[0m[38;2;29;24;21ms[0m[38;2;37;32;28mX[0m[38;2;34;26;21ms[0m[38;2;53;41;27m2[0m[38;2;78;66;47mM[0m[38;2;72;62;42mh[0m[38;2;119;109;86m9[0m[38;2;28;24;15mr[0m[38;2;23;21;17mr[0m[38;2;29;23;15mr[0m[38;2;62;47;36m5[0m[38;2;122;95;71m#[0m[38;2;180;146;108m@[0m[38;2;191;157;116m@[0m[38;2;189;156;111m@[0m[38;2;187;155;109m@[0m[38;2;187;154;111m@[0m[38;2;189;154;116m@[0m[38;2;164;131;98m&[0m[38;2;143;101;76m9[0m[38;2;157;102;81mB[0m[38;2;162;103;85mB[0m[38;2;161;105;85mB[0m[38;2;166;117;90m&[0m[38;2;182;141;105m@[0m[38;2;189;153;113m@[0m[38;2;187;153;111m@[0m[38;2;187;155;112m@[0m[38;2;188;155;113m@[0m[38;2;189;155;112m@[0m[38;2;190;154;111m@[0m[38;2;192;156;113m@[0m[38;2;191;157;113m@[0m[38;2;182;150;109m@[0m[38;2;144;116;87mB[0m[38;2;73;52;34m3[0m[38;2;99;88;67mS[0m[38;2;134;119;96mB[0m[38;2;46;39;25mA[0m[38;2;23;21;16mr[0m[38;2;27;20;17mr[0m[38;2;28;21;17mr[0m[38;2;25;22;17mr[0m[38;2;26;23;17mr[0m[38;2;27;22;17mr[0m[38;2;26;22;15mr[0m[38;2;27;23;15mr[0m[38;2;25;21;12mi[0m[38;2;38;34;23mX[0m[38;2;53;49;37m5[0m[38;2;44;38;26mA[0m[38;2;35;28;21ms[0m[38;2;22;16;12mi[0m[38;2;17;12;8m;[0m[38;2;15;12;6m:[0m[38;2;16;13;6m;[0m[38;2;16;13;6m;[0m[38;2;16;12;6m:[0m[38;2;16;13;6m;[0m[38;2;14;11;7m:[0m[38;2;28;21;13mr[0m[38;2;36;32;19mX[0m[38;2;17;9;8m:[0m[38;2;66;47;31m5[0m[38;2;161;126;93m&[0m[38;2;170;129;86m&[0m[38;2;168;130;90m&[0m[38;2;170;130;96m&[0m[38;2;153;112;87mB[0m[38;2;118;83;61mS[0m[38;2;95;66;47mH[0m[38;2;87;60;42mM[0m[38;2;83;58;36mh[0m[38;2;96;73;43mH[0m[38;2;126;98;62m#[0m[38;2;146;112;72m9[0m[38;2;149;113;71mB[0m[38;2;148;112;69m9[0m[38;2;150;112;70mB[0m[38;2;150;112;72mB[0m[38;2;149;112;73mB[0m[38;2;141;107;69m9[0m[38;2;106;76;45mG[0m[38;2;99;70;42mH[0m[38;2;106;75;47mG[0m[38;2;124;90;57m#[0m[38;2;137;99;62m#[0m[38;2;141;102;63m9[0m[38;2;140;101;61m9[0m[38;2;140;101;61m9[0m[38;2;141;100;60m9[0m[38;2;140;101;61m9[0m[38;2;138;100;60m#[0m[38;2;138;100;60m#[0m[38;2;138;100;60m#[0m[38;2;138;100;60m#[0m[38;2;138;100;61m9[0m");
	$display("[38;2;126;95;55m#[0m[38;2;127;95;56m#[0m[38;2;127;95;56m#[0m[38;2;127;95;56m#[0m[38;2;127;95;56m#[0m[38;2;127;95;56m#[0m[38;2;127;96;56m#[0m[38;2;127;95;56m#[0m[38;2;127;95;56m#[0m[38;2;128;95;56m#[0m[38;2;128;95;56m#[0m[38;2;127;95;56m#[0m[38;2;127;96;56m#[0m[38;2;127;95;56m#[0m[38;2;128;95;55m#[0m[38;2;131;97;55m#[0m[38;2;125;93;55m#[0m[38;2;108;83;52mG[0m[38;2;85;64;40mM[0m[38;2;58;40;23m2[0m[38;2;46;29;19mX[0m[38;2;58;37;28m2[0m[38;2;77;51;38mh[0m[38;2;106;76;55mG[0m[38;2;143;105;76m9[0m[38;2;160;117;87mB[0m[38;2;114;87;70m#[0m[38;2;17;9;7m:[0m[38;2;23;19;15mi[0m[38;2;35;26;19ms[0m[38;2;13;12;7m:[0m[38;2;9;10;9m:[0m[38;2;17;12;7m;[0m[38;2;23;19;12mi[0m[38;2;28;25;17mr[0m[38;2;30;27;20ms[0m[38;2;27;23;18mr[0m[38;2;21;15;10m;[0m[38;2;14;10;5m:[0m[38;2;15;12;8m;[0m[38;2;25;21;16mr[0m[38;2;20;17;14mi[0m[38;2;25;23;20mr[0m[38;2;49;41;30m2[0m[38;2;118;105;87m9[0m[38;2;31;25;18ms[0m[38;2;23;19;16mi[0m[38;2;37;32;23mX[0m[38;2;54;52;40m5[0m[38;2;21;13;6m;[0m[38;2;68;47;36m3[0m[38;2;130;103;78m9[0m[38;2;175;142;105m&[0m[38;2;193;155;112m@[0m[38;2;192;156;114m@[0m[38;2;189;155;114m@[0m[38;2;189;157;110m@[0m[38;2;191;156;111m@[0m[38;2;189;153;113m@[0m[38;2;187;154;112m@[0m[38;2;188;155;112m@[0m[38;2;191;156;114m@[0m[38;2;189;155;113m@[0m[38;2;188;155;110m@[0m[38;2;187;155;110m@[0m[38;2;188;156;110m@[0m[38;2;192;158;109m@[0m[38;2;192;157;113m@[0m[38;2;185;149;113m@[0m[38;2;165;130;98m&[0m[38;2;123;94;70m#[0m[38;2;72;50;40m3[0m[38;2;32;18;12mr[0m[38;2;42;31;18mX[0m[38;2;130;117;99mB[0m[38;2;72;65;49mM[0m[38;2;27;25;16mr[0m[38;2;22;18;14mi[0m[38;2;30;25;21ms[0m[38;2;29;26;21ms[0m[38;2;25;23;16mr[0m[38;2;26;23;15mr[0m[38;2;25;21;13mi[0m[38;2;44;36;29mA[0m[38;2;37;28;22mX[0m[38;2;34;26;18ms[0m[38;2;43;35;27mA[0m[38;2;40;34;25mX[0m[38;2;24;20;11mi[0m[38;2;15;12;5m:[0m[38;2;14;12;7m:[0m[38;2;16;13;8m;[0m[38;2;16;13;7m;[0m[38;2;16;13;6m;[0m[38;2;16;13;6m;[0m[38;2;17;12;6m;[0m[38;2;16;12;6m:[0m[38;2;16;13;5m:[0m[38;2;46;39;26mA[0m[38;2;47;38;24mA[0m[38;2;25;16;12mi[0m[38;2;32;20;11mr[0m[38;2;141;111;84mB[0m[38;2;170;130;91m&[0m[38;2;156;119;85mB[0m[38;2;120;87;62mS[0m[38;2;94;63;44mH[0m[38;2;88;61;44mM[0m[38;2;81;56;38mh[0m[38;2;92;66;43mH[0m[38;2;120;91;62m#[0m[38;2;141;108;72m9[0m[38;2;147;112;73mB[0m[38;2;146;110;70m9[0m[38;2;144;111;71m9[0m[38;2;144;112;71m9[0m[38;2;144;111;70m9[0m[38;2;144;111;70m9[0m[38;2;144;111;70m9[0m[38;2;139;107;65m9[0m[38;2;113;79;40mG[0m[38;2;122;85;49mS[0m[38;2;136;97;63m#[0m[38;2;140;101;63m9[0m[38;2;141;100;61m9[0m[38;2;141;99;59m9[0m[38;2;140;100;59m9[0m[38;2;140;100;59m9[0m[38;2;141;100;60m9[0m[38;2;141;100;60m9[0m[38;2;141;100;61m9[0m[38;2;141;100;62m9[0m[38;2;140;99;61m9[0m[38;2;139;98;60m#[0m[38;2;138;100;59m#[0m");
	$display("[38;2;125;93;54m#[0m[38;2;125;93;54m#[0m[38;2;125;93;54m#[0m[38;2;126;94;55m#[0m[38;2;126;94;55m#[0m[38;2;125;93;54m#[0m[38;2;125;93;55m#[0m[38;2;125;93;54m#[0m[38;2;125;93;54m#[0m[38;2;126;94;55m#[0m[38;2;126;94;55m#[0m[38;2;126;94;55m#[0m[38;2;126;94;55m#[0m[38;2;126;94;55m#[0m[38;2;126;93;55m#[0m[38;2;128;93;54m#[0m[38;2;126;92;55m#[0m[38;2;114;83;49mS[0m[38;2;96;68;38mH[0m[38;2;86;61;35mM[0m[38;2;70;50;28m3[0m[38;2;53;35;19mA[0m[38;2;47;30;17mX[0m[38;2;57;40;27m2[0m[38;2;79;54;35mh[0m[38;2;105;78;58mG[0m[38;2;62;46;37m5[0m[38;2;11;6;5m,[0m[38;2;33;27;19ms[0m[38;2;47;41;30m2[0m[38;2;21;20;15mi[0m[38;2;10;9;7m:[0m[38;2;12;9;8m:[0m[38;2;14;11;7m:[0m[38;2;13;11;5m:[0m[38;2;18;15;9m;[0m[38;2;24;22;17mr[0m[38;2;31;28;23ms[0m[38;2;30;27;22ms[0m[38;2;23;20;15mi[0m[38;2;15;12;7m:[0m[38;2;16;12;7m;[0m[38;2;32;29;25mX[0m[38;2;34;26;17ms[0m[38;2;107;96;78m#[0m[38;2;32;27;18ms[0m[38;2;15;14;9m;[0m[38;2;39;30;25mX[0m[38;2;60;48;43m3[0m[38;2;22;15;13mi[0m[38;2;17;13;13m;[0m[38;2;22;16;13mi[0m[38;2;46;36;28mA[0m[38;2;87;69;53mH[0m[38;2;132;105;81m9[0m[38;2;170;137;103m&[0m[38;2;187;152;107m@[0m[38;2;193;156;112m@[0m[38;2;194;156;116m@[0m[38;2;192;157;113m@[0m[38;2;191;158;113m@[0m[38;2;191;158;114m@[0m[38;2;190;157;113m@[0m[38;2;187;154;111m@[0m[38;2;180;147;106m@[0m[38;2;165;133;98m&[0m[38;2;141;111;86mB[0m[38;2;111;83;68mS[0m[38;2;78;54;43mh[0m[38;2;51;30;23mA[0m[38;2;37;19;18ms[0m[38;2;30;18;18mr[0m[38;2;29;20;12mr[0m[38;2;89;81;63mG[0m[38;2;84;74;54mH[0m[38;2;35;30;19ms[0m[38;2;18;16;11m;[0m[38;2;10;4;3m,[0m[38;2;38;29;27mX[0m[38;2;38;30;27mX[0m[38;2;25;21;15mr[0m[38;2;24;21;15mr[0m[38;2;25;21;14mr[0m[38;2;55;46;37m5[0m[38;2;50;42;33m2[0m[38;2;37;32;25mX[0m[38;2;25;22;16mr[0m[38;2;14;12;8m:[0m[38;2;14;11;7m:[0m[38;2;14;12;7m:[0m[38;2;14;12;7m:[0m[38;2;15;12;7m:[0m[38;2;15;12;7m:[0m[38;2;15;12;7m:[0m[38;2;15;12;7m:[0m[38;2;15;12;7m:[0m[38;2;15;12;8m;[0m[38;2;13;11;7m:[0m[38;2;32;28;19ms[0m[38;2;48;35;26mA[0m[38;2;40;30;23mX[0m[38;2;18;10;4m:[0m[38;2;104;81;65mS[0m[38;2;125;91;69m#[0m[38;2;81;50;32m3[0m[38;2;75;50;34m3[0m[38;2;77;54;35mh[0m[38;2;84;59;36mh[0m[38;2;113;83;55mS[0m[38;2;139;105;70m9[0m[38;2;146;109;71m9[0m[38;2;145;108;68m9[0m[38;2;145;108;69m9[0m[38;2;145;108;69m9[0m[38;2;145;107;68m9[0m[38;2;144;107;68m9[0m[38;2;144;108;68m9[0m[38;2;144;108;68m9[0m[38;2;144;108;68m9[0m[38;2;145;108;69m9[0m[38;2;143;107;67m9[0m[38;2;149;109;69m9[0m[38;2;151;109;66m9[0m[38;2;150;109;64m9[0m[38;2;149;110;64m9[0m[38;2;148;110;65m9[0m[38;2;149;110;65m9[0m[38;2;149;111;66m9[0m[38;2;149;111;66m9[0m[38;2;148;109;64m9[0m[38;2;146;108;63m9[0m[38;2;147;108;64m9[0m[38;2;146;107;64m9[0m[38;2;146;106;64m9[0m[38;2;147;106;63m9[0m");
	$display("[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;125;93;55m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;123;92;54mS[0m[38;2;123;92;54mS[0m[38;2;121;92;53mS[0m[38;2;119;87;50mS[0m[38;2;118;86;50mS[0m[38;2;113;85;49mS[0m[38;2;93;69;39mH[0m[38;2;72;51;28m3[0m[38;2;61;40;21m2[0m[38;2;55;34;18mA[0m[38;2;57;41;30m2[0m[38;2;23;16;11mi[0m[38;2;23;18;15mi[0m[38;2;46;35;28mA[0m[38;2;34;27;21ms[0m[38;2;13;13;12m;[0m[38;2;11;9;9m:[0m[38;2;12;9;9m:[0m[38;2;12;10;10m:[0m[38;2;12;11;7m:[0m[38;2;12;11;7m:[0m[38;2;12;11;9m:[0m[38;2;14;13;10m;[0m[38;2;19;18;15mi[0m[38;2;28;27;23ms[0m[38;2;28;27;22ms[0m[38;2;14;12;5m:[0m[38;2;27;25;20mr[0m[38;2;26;20;13mi[0m[38;2;80;68;54mH[0m[38;2;47;34;26mA[0m[38;2;25;12;10mi[0m[38;2;19;11;9m;[0m[38;2;37;27;26mX[0m[38;2;36;24;24ms[0m[38;2;9;6;4m,[0m[38;2;5;3;1m.[0m[38;2;1;2;2m.[0m[38;2;0;0;0m [0m[38;2;2;1;1m.[0m[38;2;34;26;21ms[0m[38;2;73;58;43mh[0m[38;2;109;87;65mS[0m[38;2;139;109;85mB[0m[38;2;150;117;87mB[0m[38;2;144;112;82mB[0m[38;2;131;101;75m9[0m[38;2;111;83;64mS[0m[38;2;89;64;51mH[0m[38;2;67;45;35m3[0m[38;2;51;30;24mA[0m[38;2;39;21;19ms[0m[38;2;35;19;18mr[0m[38;2;36;21;18ms[0m[38;2;38;23;18ms[0m[38;2;38;24;19ms[0m[38;2;32;21;17mr[0m[38;2;55;47;41m5[0m[38;2;61;55;47m3[0m[38;2;34;29;21ms[0m[38;2;19;18;14mi[0m[38;2;4;3;4m.[0m[38;2;8;5;5m,[0m[38;2;41;36;33mA[0m[38;2;34;28;25mX[0m[38;2;24;21;15mr[0m[38;2;33;32;24mX[0m[38;2;40;36;29mA[0m[38;2;32;28;21ms[0m[38;2;22;17;12mi[0m[38;2;14;11;8m:[0m[38;2;12;11;8m:[0m[38;2;12;11;10m:[0m[38;2;12;11;8m:[0m[38;2;12;11;8m:[0m[38;2;12;11;8m:[0m[38;2;12;12;7m:[0m[38;2;13;11;8m:[0m[38;2;13;11;9m:[0m[38;2;13;11;9m:[0m[38;2;13;11;8m:[0m[38;2;12;11;8m:[0m[38;2;11;11;7m:[0m[38;2;14;13;7m:[0m[38;2;45;36;28mA[0m[38;2;56;45;35m5[0m[38;2;26;22;12mr[0m[38;2;36;27;19ms[0m[38;2;52;34;25mA[0m[38;2;42;23;16ms[0m[38;2;60;36;25m2[0m[38;2;94;64;41mM[0m[38;2;126;93;64m#[0m[38;2;142;107;71m9[0m[38;2;143;107;68m9[0m[38;2;142;107;67m9[0m[38;2;142;107;68m9[0m[38;2;141;106;68m9[0m[38;2;142;106;68m9[0m[38;2;141;106;68m9[0m[38;2;141;106;67m9[0m[38;2;143;107;69m9[0m[38;2;143;107;69m9[0m[38;2;143;107;69m9[0m[38;2;143;107;69m9[0m[38;2;144;108;68m9[0m[38;2;146;109;67m9[0m[38;2;147;109;66m9[0m[38;2;145;109;65m9[0m[38;2;145;110;65m9[0m[38;2;146;109;65m9[0m[38;2;145;108;64m9[0m[38;2;145;108;64m9[0m[38;2;145;108;64m9[0m[38;2;144;107;65m9[0m[38;2;144;106;65m9[0m[38;2;143;105;65m9[0m[38;2;142;104;65m9[0m[38;2;142;104;65m9[0m[38;2;141;104;63m9[0m");
	$display("[38;2;123;91;53mS[0m[38;2;123;91;53mS[0m[38;2;123;91;53mS[0m[38;2;123;91;53mS[0m[38;2;123;91;53mS[0m[38;2;123;91;53mS[0m[38;2;123;91;53mS[0m[38;2;124;91;53mS[0m[38;2;124;92;54m#[0m[38;2;122;92;54mS[0m[38;2;122;92;54mS[0m[38;2;122;92;54mS[0m[38;2;122;92;54mS[0m[38;2;121;91;53mS[0m[38;2;121;91;53mS[0m[38;2;121;91;53mS[0m[38;2;120;91;53mS[0m[38;2;121;91;53mS[0m[38;2;122;91;54mS[0m[38;2;123;92;53mS[0m[38;2;117;88;50mS[0m[38;2;97;72;39mH[0m[38;2;87;63;37mM[0m[38;2;96;71;47mH[0m[38;2;80;55;32mh[0m[38;2;52;36;23mA[0m[38;2;17;12;5m:[0m[38;2;45;38;26mA[0m[38;2;61;49;35m5[0m[38;2;31;26;18ms[0m[38;2;12;11;8m:[0m[38;2;12;11;7m:[0m[38;2;10;11;8m:[0m[38;2;11;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;8m:[0m[38;2;11;12;7m:[0m[38;2;12;11;8m:[0m[38;2;12;11;9m:[0m[38;2;14;13;10m;[0m[38;2;20;19;14mi[0m[38;2;18;18;10m;[0m[38;2;22;22;17mr[0m[38;2;26;24;20mr[0m[38;2;39;30;24mX[0m[38;2;63;46;36m5[0m[38;2;105;67;59mG[0m[38;2;60;23;22mA[0m[38;2;18;10;9m;[0m[38;2;11;5;6m,[0m[38;2;4;4;3m.[0m[38;2;0;1;1m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;1m.[0m[38;2;0;1;2m.[0m[38;2;12;11;9m:[0m[38;2;21;15;9m;[0m[38;2;28;16;12mi[0m[38;2;39;23;23ms[0m[38;2;38;22;20ms[0m[38;2;38;19;18ms[0m[38;2;37;18;17mr[0m[38;2;35;20;17mr[0m[38;2;34;22;19ms[0m[38;2;37;23;21ms[0m[38;2;38;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;38;23;21ms[0m[38;2;34;22;19ms[0m[38;2;30;21;17mr[0m[38;2;31;26;21ms[0m[38;2;27;24;18mr[0m[38;2;17;16;12m;[0m[38;2;4;3;2m.[0m[38;2;1;0;0m.[0m[38;2;5;4;3m,[0m[38;2;16;14;13m;[0m[38;2;14;9;8m:[0m[38;2;29;27;21ms[0m[38;2;38;40;30mA[0m[38;2;23;18;11mi[0m[38;2;13;9;7m:[0m[38;2;13;9;8m:[0m[38;2;13;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;8m:[0m[38;2;12;11;7m:[0m[38;2;50;40;29m2[0m[38;2;76;61;44mh[0m[38;2;38;30;18mX[0m[38;2;20;13;12m;[0m[38;2;34;24;17ms[0m[38;2;20;8;6m:[0m[38;2;60;39;30m2[0m[38;2;117;82;59mS[0m[38;2;133;97;67m#[0m[38;2;139;105;67m9[0m[38;2;139;106;65m9[0m[38;2;138;105;65m9[0m[38;2;139;105;67m9[0m[38;2;140;106;68m9[0m[38;2;139;106;68m9[0m[38;2;138;104;66m9[0m[38;2;139;104;66m9[0m[38;2;139;104;66m9[0m[38;2;140;105;67m9[0m[38;2;139;105;67m9[0m[38;2;139;104;66m9[0m[38;2;141;104;66m9[0m[38;2;143;106;65m9[0m[38;2;143;106;63m9[0m[38;2;144;107;65m9[0m[38;2;144;107;65m9[0m[38;2;143;106;64m9[0m[38;2;143;106;64m9[0m[38;2;143;106;63m9[0m[38;2;142;105;62m9[0m[38;2;142;104;65m9[0m[38;2;142;104;65m9[0m[38;2;141;103;64m9[0m[38;2;139;101;62m9[0m[38;2;140;102;63m9[0m[38;2;140;102;63m9[0m");
	$display("[38;2;122;89;52mS[0m[38;2;122;90;52mS[0m[38;2;122;90;52mS[0m[38;2;122;89;52mS[0m[38;2;121;89;52mS[0m[38;2;120;89;52mS[0m[38;2;120;90;52mS[0m[38;2;121;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;121;90;53mS[0m[38;2;122;90;52mS[0m[38;2;116;89;51mS[0m[38;2;99;74;41mH[0m[38;2;85;61;35mh[0m[38;2;96;71;45mH[0m[38;2;95;69;40mH[0m[38;2;76;59;38mh[0m[38;2;28;20;8mi[0m[38;2;60;51;36m3[0m[38;2;79;66;47mM[0m[38;2;44;35;25mA[0m[38;2;23;19;13mi[0m[38;2;17;17;11m;[0m[38;2;14;16;10m;[0m[38;2;16;16;12m;[0m[38;2;18;16;11m;[0m[38;2;19;17;11mi[0m[38;2;17;17;10m;[0m[38;2;14;14;8m;[0m[38;2;13;12;8m:[0m[38;2;12;11;8m:[0m[38;2;13;13;8m:[0m[38;2;20;17;11mi[0m[38;2;24;16;11mi[0m[38;2;39;31;24mX[0m[38;2;49;41;31m2[0m[38;2;31;21;9mr[0m[38;2;58;14;13ms[0m[38;2;58;3;9mr[0m[38;2;13;1;0m,[0m[38;2;4;4;3m.[0m[38;2;11;11;12m:[0m[38;2;8;8;8m:[0m[38;2;2;2;2m.[0m[38;2;1;1;1m.[0m[38;2;1;1;1m.[0m[38;2;0;1;0m.[0m[38;2;2;2;1m.[0m[38;2;16;12;9m;[0m[38;2;27;17;15mi[0m[38;2;36;23;23ms[0m[38;2;36;24;21ms[0m[38;2;38;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;24;20ms[0m[38;2;39;24;20ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;37;22;19ms[0m[38;2;35;22;20ms[0m[38;2;30;20;19mr[0m[38;2;24;18;16mi[0m[38;2;21;17;14mi[0m[38;2;5;4;1m.[0m[38;2;1;0;0m.[0m[38;2;6;4;5m,[0m[38;2;12;11;10m:[0m[38;2;10;8;8m:[0m[38;2;8;8;6m,[0m[38;2;15;13;9m;[0m[38;2;23;16;13mi[0m[38;2;12;10;7m:[0m[38;2;14;10;9m:[0m[38;2;14;10;9m:[0m[38;2;13;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;8m:[0m[38;2;12;11;8m:[0m[38;2;11;11;7m:[0m[38;2;34;26;17ms[0m[38;2;49;37;24mA[0m[38;2;32;26;16ms[0m[38;2;14;8;11m:[0m[38;2;10;6;4m,[0m[38;2;5;0;0m.[0m[38;2;60;43;32m5[0m[38;2;113;79;54mS[0m[38;2;130;94;63m#[0m[38;2;136;102;65m9[0m[38;2;137;104;65m9[0m[38;2;136;102;65m9[0m[38;2;136;102;64m9[0m[38;2;135;101;63m9[0m[38;2;135;101;63m9[0m[38;2;135;101;64m9[0m[38;2;135;101;63m9[0m[38;2;135;101;63m9[0m[38;2;136;101;63m9[0m[38;2;136;102;64m9[0m[38;2;137;103;65m9[0m[38;2;139;102;65m9[0m[38;2;140;104;63m9[0m[38;2;140;104;61m9[0m[38;2;140;104;62m9[0m[38;2;141;104;64m9[0m[38;2;141;103;63m9[0m[38;2;140;103;62m9[0m[38;2;140;103;62m9[0m[38;2;139;102;61m9[0m[38;2;139;101;62m9[0m[38;2;139;101;62m9[0m[38;2;138;100;61m9[0m[38;2;136;98;59m#[0m[38;2;138;99;60m#[0m[38;2;139;101;62m9[0m");
	$display("[38;2;119;89;50mS[0m[38;2;119;89;49mS[0m[38;2;119;89;49mS[0m[38;2;119;89;50mS[0m[38;2;118;89;50mS[0m[38;2;118;89;50mS[0m[38;2;118;89;49mS[0m[38;2;118;89;50mS[0m[38;2;119;89;50mS[0m[38;2;120;89;50mS[0m[38;2;120;89;50mS[0m[38;2;120;89;50mS[0m[38;2;120;89;50mS[0m[38;2;120;89;50mS[0m[38;2;119;89;50mS[0m[38;2;118;89;49mS[0m[38;2;118;89;50mS[0m[38;2;118;89;49mS[0m[38;2;118;88;51mS[0m[38;2;119;88;50mS[0m[38;2;118;87;50mS[0m[38;2;103;77;45mG[0m[38;2;84;62;36mM[0m[38;2;92;68;41mH[0m[38;2;87;61;33mh[0m[38;2;71;53;32m3[0m[38;2;44;32;21mX[0m[38;2;57;47;35m5[0m[38;2;57;46;31m5[0m[38;2;47;36;26mA[0m[38;2;40;32;25mX[0m[38;2;29;25;18mr[0m[38;2;25;24;17mr[0m[38;2;28;25;19mr[0m[38;2;34;28;21ms[0m[38;2;37;30;22mX[0m[38;2;38;33;24mX[0m[38;2;36;31;24mX[0m[38;2;29;23;19mr[0m[38;2;19;15;12m;[0m[38;2;20;14;11m;[0m[38;2;35;9;7mi[0m[38;2;64;29;24m2[0m[38;2;55;28;21mA[0m[38;2;57;27;21mA[0m[38;2;40;13;8mr[0m[38;2;44;12;12mr[0m[38;2;59;7;15ms[0m[38;2;34;5;8mi[0m[38;2;12;9;6m:[0m[38;2;12;9;8m:[0m[38;2;10;10;9m:[0m[38;2;3;3;2m.[0m[38;2;1;1;1m.[0m[38;2;1;1;1m.[0m[38;2;1;1;1m.[0m[38;2;1;0;1m.[0m[38;2;5;0;1m.[0m[38;2;26;15;14mi[0m[38;2;39;22;20ms[0m[38;2;37;22;18ms[0m[38;2;37;23;19ms[0m[38;2;38;23;20ms[0m[38;2;39;22;20ms[0m[38;2;39;22;20ms[0m[38;2;38;23;20ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;23;22ms[0m[38;2;36;22;21ms[0m[38;2;22;15;13mi[0m[38;2;8;7;5m,[0m[38;2;4;3;3m.[0m[38;2;11;10;10m:[0m[38;2;18;16;16mi[0m[38;2;15;12;12m;[0m[38;2;4;2;1m.[0m[38;2;1;3;1m.[0m[38;2;19;4;3m:[0m[38;2;38;4;7mi[0m[38;2;19;9;9m;[0m[38;2;11;12;8m:[0m[38;2;13;11;8m:[0m[38;2;12;11;8m:[0m[38;2;12;11;9m:[0m[38;2;14;10;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;12;10;8m:[0m[38;2;15;11;3m:[0m[38;2;31;28;20ms[0m[38;2;23;22;18mr[0m[38;2;10;7;8m:[0m[38;2;4;1;2m.[0m[38;2;8;1;1m.[0m[38;2;67;47;36m3[0m[38;2;108;76;49mG[0m[38;2;126;92;57m#[0m[38;2;134;98;63m#[0m[38;2;136;100;66m9[0m[38;2;133;99;62m#[0m[38;2;132;98;60m#[0m[38;2;132;98;60m#[0m[38;2;132;98;61m#[0m[38;2;132;98;61m#[0m[38;2;132;98;60m#[0m[38;2;133;99;62m#[0m[38;2;134;100;62m#[0m[38;2;134;100;62m#[0m[38;2;134;100;62m#[0m[38;2;135;100;63m#[0m[38;2;137;102;64m9[0m[38;2;137;102;64m9[0m[38;2;137;102;64m9[0m[38;2;137;102;64m9[0m[38;2;137;101;64m9[0m[38;2;137;100;63m9[0m[38;2;138;99;63m9[0m[38;2;137;99;62m#[0m[38;2;137;99;61m#[0m[38;2;137;98;61m#[0m[38;2;137;99;61m#[0m[38;2;137;98;59m#[0m[38;2;137;98;59m#[0m[38;2;137;98;59m#[0m");
	$display("[38;2;117;88;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;49mS[0m[38;2;117;88;49mS[0m[38;2;117;87;49mS[0m[38;2;118;88;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;49mS[0m[38;2;118;87;49mS[0m[38;2;118;87;49mS[0m[38;2;118;87;49mS[0m[38;2;118;88;49mS[0m[38;2;118;87;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;50mS[0m[38;2;118;87;49mS[0m[38;2;118;86;49mS[0m[38;2;105;79;46mG[0m[38;2;86;65;39mM[0m[38;2;90;67;42mM[0m[38;2;84;57;31mh[0m[38;2;75;56;36mh[0m[38;2;44;34;23mA[0m[38;2;45;36;25mA[0m[38;2;52;43;29m2[0m[38;2;51;41;30m2[0m[38;2;35;27;18ms[0m[38;2;27;24;17mr[0m[38;2;24;21;15mr[0m[38;2;25;20;15mr[0m[38;2;29;21;17mr[0m[38;2;31;23;20ms[0m[38;2;32;25;20ms[0m[38;2;33;25;21ms[0m[38;2;28;24;21ms[0m[38;2;23;18;14mi[0m[38;2;39;8;8mi[0m[38;2;71;21;17mA[0m[38;2;137;94;80m9[0m[38;2;65;30;20m2[0m[38;2;53;10;8mr[0m[38;2;62;8;12ms[0m[38;2;48;9;13mr[0m[38;2;30;9;11mi[0m[38;2;15;10;10m;[0m[38;2;10;10;10m:[0m[38;2;11;9;9m:[0m[38;2;11;11;9m:[0m[38;2;4;4;3m.[0m[38;2;1;1;1m.[0m[38;2;1;1;1m.[0m[38;2;1;1;1m.[0m[38;2;2;1;1m.[0m[38;2;4;0;1m.[0m[38;2;26;14;14mi[0m[38;2;38;20;19ms[0m[38;2;35;19;16mr[0m[38;2;35;20;17mr[0m[38;2;35;19;17mr[0m[38;2;36;20;19ms[0m[38;2;36;20;19ms[0m[38;2;37;22;20ms[0m[38;2;37;22;19ms[0m[38;2;37;22;19ms[0m[38;2;37;22;19ms[0m[38;2;38;22;21ms[0m[38;2;40;23;23mX[0m[38;2;29;15;15mi[0m[38;2;10;3;2m,[0m[38;2;10;9;6m:[0m[38;2;13;15;10m;[0m[38;2;13;13;9m;[0m[38;2;13;10;7m:[0m[38;2;14;8;6m:[0m[38;2;18;3;5m:[0m[38;2;31;7;7m;[0m[38;2;105;67;57mG[0m[38;2;91;41;32mh[0m[38;2;45;2;5mi[0m[38;2;19;9;6m:[0m[38;2;10;11;6m:[0m[38;2;12;10;9m:[0m[38;2;12;9;9m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;10;10;8m:[0m[38;2;16;11;11m;[0m[38;2;44;39;30mA[0m[38;2;35;30;21mX[0m[38;2;14;11;9m:[0m[38;2;11;6;6m:[0m[38;2;4;0;1m.[0m[38;2;11;4;2m,[0m[38;2;74;55;40mh[0m[38;2;106;75;46mG[0m[38;2;123;90;53mS[0m[38;2;132;97;60m#[0m[38;2;132;97;62m#[0m[38;2;130;97;59m#[0m[38;2;129;95;58m#[0m[38;2;129;95;58m#[0m[38;2;131;97;60m#[0m[38;2;130;96;59m#[0m[38;2;130;96;59m#[0m[38;2;131;97;60m#[0m[38;2;130;96;59m#[0m[38;2;131;97;59m#[0m[38;2;132;98;60m#[0m[38;2;133;99;61m#[0m[38;2;134;100;62m#[0m[38;2;134;100;62m#[0m[38;2;134;99;61m#[0m[38;2;134;99;61m#[0m[38;2;134;99;61m#[0m[38;2;135;98;61m#[0m[38;2;136;98;61m#[0m[38;2;135;97;60m#[0m[38;2;134;98;60m#[0m[38;2;134;98;61m#[0m[38;2;135;99;60m#[0m[38;2;133;98;58m#[0m[38;2;133;97;58m#[0m[38;2;133;97;58m#[0m");
	$display("[38;2;115;85;49mS[0m[38;2;116;86;49mS[0m[38;2;116;86;49mS[0m[38;2;115;85;49mS[0m[38;2;115;85;49mS[0m[38;2;115;86;49mS[0m[38;2;116;87;50mS[0m[38;2;116;86;50mS[0m[38;2;116;86;50mS[0m[38;2;115;87;50mS[0m[38;2;115;87;50mS[0m[38;2;115;87;50mS[0m[38;2;115;87;50mS[0m[38;2;116;87;50mS[0m[38;2;116;86;50mS[0m[38;2;116;86;50mS[0m[38;2;116;86;50mS[0m[38;2;116;86;50mS[0m[38;2;116;86;50mS[0m[38;2;117;86;48mS[0m[38;2;116;85;48mS[0m[38;2;107;80;48mG[0m[38;2;89;67;41mM[0m[38;2;89;67;44mM[0m[38;2;82;55;29mh[0m[38;2;83;62;41mM[0m[38;2;30;23;11mr[0m[38;2;26;22;14mr[0m[38;2;47;38;28mA[0m[38;2;47;38;31m2[0m[38;2;18;11;8m;[0m[38;2;14;11;9m:[0m[38;2;12;11;8m:[0m[38;2;11;10;7m:[0m[38;2;12;9;7m:[0m[38;2;10;9;8m:[0m[38;2;9;9;7m:[0m[38;2;10;8;6m:[0m[38;2;11;9;10m:[0m[38;2;20;6;7m:[0m[38;2;49;5;4mi[0m[38;2;131;76;65m#[0m[38;2;124;69;58mS[0m[38;2;70;6;8ms[0m[38;2;65;5;9ms[0m[38;2;66;3;8ms[0m[38;2;49;4;7mr[0m[38;2;9;4;2m,[0m[38;2;5;8;7m,[0m[38;2;13;7;7m:[0m[38;2;9;9;6m:[0m[38;2;10;10;8m:[0m[38;2;7;7;5m,[0m[38;2;0;1;0m.[0m[38;2;1;1;1m.[0m[38;2;1;2;1m.[0m[38;2;1;1;2m.[0m[38;2;4;0;0m.[0m[38;2;46;31;28mA[0m[38;2;62;41;34m5[0m[38;2;82;61;47mM[0m[38;2;78;58;43mh[0m[38;2;85;66;53mH[0m[38;2;61;42;32m5[0m[38;2;57;39;31m2[0m[38;2;38;21;18ms[0m[38;2;37;21;19ms[0m[38;2;38;22;20ms[0m[38;2;37;23;20ms[0m[38;2;32;21;20ms[0m[38;2;23;14;13mi[0m[38;2;9;3;2m,[0m[38;2;9;6;5m,[0m[38;2;12;10;9m:[0m[38;2;12;9;8m:[0m[38;2;12;9;9m:[0m[38;2;13;9;9m:[0m[38;2;13;9;10m:[0m[38;2;20;6;5m:[0m[38;2;41;1;2m;[0m[38;2;86;38;34m3[0m[38;2;145;102;87mB[0m[38;2;84;28;23m5[0m[38;2;43;3;4mi[0m[38;2;14;9;6m:[0m[38;2;7;11;10m:[0m[38;2;13;8;10m:[0m[38;2;12;9;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;10;9;7m:[0m[38;2;16;12;11m;[0m[38;2;41;33;26mA[0m[38;2;43;34;27mA[0m[38;2;18;14;12m;[0m[38;2;9;7;6m,[0m[38;2;4;0;0m.[0m[38;2;21;11;7m;[0m[38;2;84;59;42mM[0m[38;2;101;71;43mH[0m[38;2;120;88;53mS[0m[38;2;128;95;59m#[0m[38;2;129;95;61m#[0m[38;2;127;95;58m#[0m[38;2;127;93;57m#[0m[38;2;127;93;57m#[0m[38;2;128;94;58m#[0m[38;2;126;92;57m#[0m[38;2;127;93;56m#[0m[38;2;128;94;57m#[0m[38;2;128;94;56m#[0m[38;2;129;95;57m#[0m[38;2;129;95;57m#[0m[38;2;129;95;58m#[0m[38;2;131;97;60m#[0m[38;2;130;96;59m#[0m[38;2;130;96;59m#[0m[38;2;131;96;59m#[0m[38;2;133;97;59m#[0m[38;2;134;97;60m#[0m[38;2;135;97;60m#[0m[38;2;135;96;59m#[0m[38;2;134;96;59m#[0m[38;2;133;95;58m#[0m[38;2;133;95;57m#[0m[38;2;131;94;55m#[0m[38;2;130;93;55m#[0m[38;2;130;94;56m#[0m");
	$display("[38;2;115;85;49mS[0m[38;2;115;85;49mS[0m[38;2;114;84;48mS[0m[38;2;115;85;49mS[0m[38;2;115;85;49mS[0m[38;2;114;86;49mS[0m[38;2;115;87;50mS[0m[38;2;114;86;49mS[0m[38;2;114;86;49mS[0m[38;2;114;86;49mS[0m[38;2;115;87;50mS[0m[38;2;115;87;50mS[0m[38;2;114;86;49mS[0m[38;2;114;86;49mS[0m[38;2;115;85;49mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;109;81;50mG[0m[38;2;93;69;41mH[0m[38;2;84;61;36mh[0m[38;2;81;56;27mh[0m[38;2;94;73;47mH[0m[38;2;33;23;12mr[0m[38;2;23;18;14mi[0m[38;2;55;44;32m5[0m[38;2;43;34;24mA[0m[38;2;15;9;8m:[0m[38;2;11;8;8m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;9;9;7m:[0m[38;2;16;5;9m:[0m[38;2;35;2;6m;[0m[38;2;83;36;30m3[0m[38;2;151;100;85mB[0m[38;2;82;21;17m2[0m[38;2;71;4;9ms[0m[38;2;69;2;5ms[0m[38;2;66;2;5ms[0m[38;2;52;3;5mr[0m[38;2;16;2;3m,[0m[38;2;6;6;7m,[0m[38;2;15;10;9m:[0m[38;2;19;15;15mi[0m[38;2;18;15;13m;[0m[38;2;14;14;10m;[0m[38;2;7;6;3m,[0m[38;2;5;2;3m.[0m[38;2;1;1;3m.[0m[38;2;1;1;1m.[0m[38;2;53;39;31m2[0m[38;2;128;105;86m9[0m[38;2;100;81;61mG[0m[38;2;105;86;67mS[0m[38;2;108;85;68mS[0m[38;2;110;85;67mS[0m[38;2;132;108;83m9[0m[38;2;146;119;94mB[0m[38;2;81;57;45mM[0m[38;2;34;18;15mr[0m[38;2;30;17;16mr[0m[38;2;20;14;11m;[0m[38;2;8;7;4m,[0m[38;2;6;5;2m,[0m[38;2;9;7;6m,[0m[38;2;11;9;8m:[0m[38;2;11;10;9m:[0m[38;2;12;10;8m:[0m[38;2;11;10;8m:[0m[38;2;10;10;8m:[0m[38;2;7;8;6m,[0m[38;2;15;5;3m:[0m[38;2;42;3;4mi[0m[38;2;51;0;0mi[0m[38;2;106;60;51mH[0m[38;2;141;96;79m9[0m[38;2;62;13;11mX[0m[38;2;30;5;3m;[0m[38;2;10;9;5m:[0m[38;2;10;10;7m:[0m[38;2;12;9;7m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;10;9;7m:[0m[38;2;15;11;8m:[0m[38;2;46;32;24mA[0m[38;2;54;41;30m2[0m[38;2;24;19;12mi[0m[38;2;6;5;4m,[0m[38;2;3;0;1m.[0m[38;2;35;21;16mr[0m[38;2;85;59;41mM[0m[38;2;99;69;42mH[0m[38;2;116;84;54mS[0m[38;2;124;91;57m#[0m[38;2;125;93;57m#[0m[38;2;123;92;56m#[0m[38;2;124;90;55mS[0m[38;2;124;90;55mS[0m[38;2;124;90;55mS[0m[38;2;124;90;55mS[0m[38;2;125;91;56m#[0m[38;2;125;91;56m#[0m[38;2;125;91;55m#[0m[38;2;125;91;54m#[0m[38;2;126;92;55m#[0m[38;2;126;92;55m#[0m[38;2;127;93;56m#[0m[38;2;127;93;56m#[0m[38;2;127;93;56m#[0m[38;2;127;93;56m#[0m[38;2;129;93;57m#[0m[38;2;129;94;56m#[0m[38;2;129;94;56m#[0m[38;2;129;93;56m#[0m[38;2;129;93;56m#[0m[38;2;129;93;56m#[0m[38;2;129;93;56m#[0m[38;2;128;92;55m#[0m[38;2;127;91;54m#[0m[38;2;127;92;54m#[0m");
	$display("[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;85;48mS[0m[38;2;114;86;48mS[0m[38;2;114;86;49mS[0m[38;2;114;86;49mS[0m[38;2;114;86;49mS[0m[38;2;114;85;49mS[0m[38;2;115;86;49mS[0m[38;2;114;85;49mS[0m[38;2;113;84;48mS[0m[38;2;113;84;48mS[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;48mG[0m[38;2;110;83;51mG[0m[38;2;95;71;43mH[0m[38;2;79;58;32mh[0m[38;2;88;61;29mh[0m[38;2;107;80;50mG[0m[38;2;54;40;26m2[0m[38;2;18;12;10m;[0m[38;2;57;47;37m5[0m[38;2;57;51;38m5[0m[38;2;19;16;11m;[0m[38;2;9;8;6m:[0m[38;2;9;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;12;8;8m:[0m[38;2;23;2;3m:[0m[38;2;47;3;3mi[0m[38;2;126;80;71m#[0m[38;2;114;66;56mG[0m[38;2;61;1;1mr[0m[38;2;62;2;5mr[0m[38;2;61;1;2mr[0m[38;2;60;0;5mr[0m[38;2;54;1;5mr[0m[38;2;38;2;8mi[0m[38;2;17;2;4m:[0m[38;2;12;7;5m:[0m[38;2;14;10;10m:[0m[38;2;15;12;9m;[0m[38;2;14;13;8m;[0m[38;2;14;13;8m;[0m[38;2;14;11;10m;[0m[38;2;11;8;9m:[0m[38;2;12;7;5m:[0m[38;2;87;72;61mH[0m[38;2;84;69;52mH[0m[38;2;42;39;24mA[0m[38;2;40;49;32m2[0m[38;2;38;43;23mA[0m[38;2;86;67;49mH[0m[38;2;149;120;98mB[0m[38;2;126;104;82m9[0m[38;2;64;51;41m3[0m[38;2;20;16;13mi[0m[38;2;17;13;10m;[0m[38;2;12;9;5m:[0m[38;2;12;11;7m:[0m[38;2;14;13;10m;[0m[38;2;16;15;13m;[0m[38;2;17;15;13m;[0m[38;2;21;19;18mi[0m[38;2;23;21;20mr[0m[38;2;23;21;18mr[0m[38;2;22;16;14mi[0m[38;2;19;6;6m:[0m[38;2;31;2;4m;[0m[38;2;49;3;8mr[0m[38;2;56;0;3mi[0m[38;2;60;6;3mr[0m[38;2;133;91;78m9[0m[38;2;114;65;56mG[0m[38;2;49;2;2mi[0m[38;2;24;5;5m:[0m[38;2;9;10;7m:[0m[38;2;10;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;10;9;7m:[0m[38;2;26;23;16mr[0m[38;2;67;55;39m3[0m[38;2;60;48;32m5[0m[38;2;19;14;7m;[0m[38;2;4;3;2m.[0m[38;2;5;1;2m.[0m[38;2;46;33;24mA[0m[38;2;82;58;36mh[0m[38;2;96;67;37mM[0m[38;2;112;80;48mG[0m[38;2;122;88;54mS[0m[38;2;123;90;56mS[0m[38;2;120;88;55mS[0m[38;2;122;87;53mS[0m[38;2;122;87;53mS[0m[38;2;122;87;53mS[0m[38;2;121;86;53mS[0m[38;2;121;87;52mS[0m[38;2;122;88;53mS[0m[38;2;122;88;52mS[0m[38;2;123;88;51mS[0m[38;2;123;89;52mS[0m[38;2;124;89;53mS[0m[38;2;126;90;54m#[0m[38;2;125;90;53mS[0m[38;2;126;90;54m#[0m[38;2;126;91;54m#[0m[38;2;126;91;54m#[0m[38;2;126;91;54m#[0m[38;2;126;92;54m#[0m[38;2;126;92;54m#[0m[38;2;126;92;54m#[0m[38;2;126;91;54m#[0m[38;2;126;91;54m#[0m[38;2;125;90;53mS[0m[38;2;124;89;52mS[0m[38;2;125;89;52mS[0m");
	$display("[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;46mG[0m[38;2;112;84;47mG[0m[38;2;111;84;48mG[0m[38;2;112;83;48mG[0m[38;2;112;83;47mG[0m[38;2;112;84;47mG[0m[38;2;112;84;47mG[0m[38;2;112;84;47mG[0m[38;2;112;84;47mG[0m[38;2;112;83;47mG[0m[38;2;111;82;46mG[0m[38;2;111;82;46mG[0m[38;2;111;82;46mG[0m[38;2;112;82;46mG[0m[38;2;112;82;46mG[0m[38;2;111;82;49mG[0m[38;2;107;82;51mG[0m[38;2;95;72;42mH[0m[38;2;79;59;29mh[0m[38;2;90;65;37mM[0m[38;2;108;79;49mG[0m[38;2;83;64;43mM[0m[38;2;17;10;6m:[0m[38;2;30;23;20ms[0m[38;2;31;26;19ms[0m[38;2;13;11;5m:[0m[38;2;9;8;4m,[0m[38;2;9;8;5m,[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;14;7;7m:[0m[38;2;30;2;1m:[0m[38;2;64;20;17mA[0m[38;2;143;98;88m9[0m[38;2;78;29;23m5[0m[38;2;55;0;2mi[0m[38;2;56;0;4mr[0m[38;2;54;1;3mi[0m[38;2;51;1;4mi[0m[38;2;49;1;1mi[0m[38;2;48;2;4mi[0m[38;2;40;2;4m;[0m[38;2;20;2;1m:[0m[38;2;6;5;3m,[0m[38;2;5;7;4m,[0m[38;2;7;8;6m,[0m[38;2;12;10;10m:[0m[38;2;14;10;9m:[0m[38;2;15;9;9m:[0m[38;2;14;10;9m:[0m[38;2;36;29;24mX[0m[38;2;46;40;28mA[0m[38;2;31;34;24mX[0m[38;2;24;34;19ms[0m[38;2;40;46;27mA[0m[38;2;69;56;41mh[0m[38;2;77;60;49mM[0m[38;2;39;30;24mX[0m[38;2;7;3;3m,[0m[38;2;9;10;9m:[0m[38;2;11;10;8m:[0m[38;2;14;11;8m:[0m[38;2;17;13;10m;[0m[38;2;15;11;8m:[0m[38;2;13;9;7m:[0m[38;2;12;8;7m:[0m[38;2;12;9;7m:[0m[38;2;12;8;6m:[0m[38;2;18;3;3m:[0m[38;2;31;1;3m;[0m[38;2;44;3;5mi[0m[38;2;49;2;4mi[0m[38;2;53;1;4mi[0m[38;2;56;0;6mr[0m[38;2;53;0;0mi[0m[38;2;88;39;36m3[0m[38;2;145;103;88mB[0m[38;2;68;19;16mA[0m[38;2;31;2;5m;[0m[38;2;11;7;8m:[0m[38;2;9;9;9m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;9;8;7m:[0m[38;2;10;9;6m:[0m[38;2;10;9;5m:[0m[38;2;10;9;5m:[0m[38;2;10;8;5m:[0m[38;2;19;15;11m;[0m[38;2;41;35;25mA[0m[38;2;30;25;17mr[0m[38;2;10;6;6m,[0m[38;2;4;1;2m.[0m[38;2;15;10;6m:[0m[38;2;58;42;26m2[0m[38;2;79;59;31mh[0m[38;2;91;66;36mM[0m[38;2;106;77;46mG[0m[38;2;114;84;51mS[0m[38;2;115;85;52mS[0m[38;2;112;82;52mS[0m[38;2;113;81;51mS[0m[38;2;112;82;51mS[0m[38;2;111;82;51mG[0m[38;2;111;81;50mG[0m[38;2;111;81;48mG[0m[38;2;113;82;49mG[0m[38;2;115;83;49mS[0m[38;2;114;83;49mS[0m[38;2;113;83;49mS[0m[38;2;114;83;48mS[0m[38;2;116;84;50mS[0m[38;2;116;85;50mS[0m[38;2;115;84;49mS[0m[38;2;115;84;49mS[0m[38;2;115;84;49mS[0m[38;2;115;84;49mS[0m[38;2;115;84;49mS[0m[38;2;115;84;49mS[0m[38;2;115;83;49mS[0m[38;2;115;84;49mS[0m[38;2;115;83;49mS[0m[38;2;115;83;48mS[0m[38;2;115;82;48mS[0m[38;2;114;82;48mG[0m");
	$display("\033[0;32m \033[5m    //   ) )     // | |     //   ) )     //   ) )\033[m");
    $display("\033[0;32m \033[5m   //___/ /     //__| |    ((           ((\033[m");
    $display("\033[0;32m \033[5m  / ____ /     / ___  |      \\           \\\033[m");
    $display("\033[0;32m \033[5m //           //    | |        ) )          ) )\033[m");
    $display("\033[0;32m \033[5m//           //     | | ((___ / /    ((___ / /\033[m");
	$display("**************************************************");
	$display("                  Congratulations!                ");
	$display("              execution cycles = %7d", total_latency);
	$display("              clock period = %4fns", CYCLE);
	$display("**************************************************");
end endtask
IFFT256 ifft_256(
    .clk(clk),
    .rst_n(rst_n),
    .in_valid(in_valid),
    .x_real(in_xp_real),
    .x_img(in_xp_img),
    .y_real(out_yp_real),
    .y_img(out_yp_img),
    .out_valid(out_valid)
);
endmodule

/*
task cal_gold_task;
    integer N;
    real    PI;
    real    scale;

    real xr [0:255];
    real xi [0:255];

    integer n, k;
    real    sumr, sumi;
    real    angle, c, s;

    integer tmp_r, tmp_i;

begin
    N     = 256;
    PI    = 3.141592653589793;
    scale = 1.0 / 256.0;

    // 1) Q1.15 array -> real
    for (n = 0; n < N; n = n + 1) begin
        xr[n] = $itor(xp_real_reg[n]) / 32768.0;  
        xi[n] = $itor(xp_img_reg[n])  / 32768.0;  
    end

    // ================================================
    // 2) 用 DFT 公式算 256 點 FFT
    //    Y[k] = Σ x[n] * exp(-j*2πkn/N)
    // ================================================
    for (k = 0; k < N; k = k + 1) begin
        sumr = 0.0;
        sumi = 0.0;

        for (n = 0; n < N; n = n + 1) begin
            angle = -2.0 * PI * $itor(k) * $itor(n) / $itor(N);
            c     = $cos(angle);
            s     = $sin(angle);

            // (xr + j*xi) * (c + j*s)
            sumr = sumr + (xr[n]*c - xi[n]*s);
            sumi = sumi + (xr[n]*s + xi[n]*c);
        end

        // 硬體如果有總體 /256，就在這裡 scale
        sumr = sumr * scale;
        sumi = sumi * scale;

        // ============================================
        // 3) real -> Q1.15，直接寫到 golden 陣列
        // ============================================
        tmp_r = $rtoi(sumr * 32768.0);  // * 2^15
        tmp_i = $rtoi(sumi * 32768.0);

        // saturation 到 Q1.15 範圍
        if (tmp_r >  32767) tmp_r =  32767;
        if (tmp_r < -32768) tmp_r = -32768;
        if (tmp_i >  32767) tmp_i =  32767;
        if (tmp_i < -32768) tmp_i = -32768;

        golden_out_yp_real[k] = tmp_r[15:0];
        golden_out_yp_img[k]  = tmp_i[15:0];
    end
end
endtask
*/